��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C���7j���Eb�Q��gQ� Q ��������˻X�"��ű��\t"�s;�K:��L%�$�������o6��)H���о��8��1c����I�#}�LB�F�P��F�r�R����]��)+?kp[�}�,:n�[�h��ٍ(>a����[��h���ߨ�I-�OeY&fދG������~��1S�S�Qi���w-�Ic��(�d��rc�3p
�-��D��!Y�L� �.��.��$�W9vCg��,\��(ݫ�2fӢ~�T&-^��A���#֩W�l9��8��Nʷ�zgy�"7����x� �]�}�MV��&Ae~�!��Z]�	<���t6hΧ̠k�m�9�c(�M;����K3����4:n(S��d�����|�5�k#��4׸�ʯ9n��r]��)s�b&&�UF�n|�'���Fz��Ɖ�a3?~ȅT�?�e�0��?��̿�{���3������* �v}5�� �Ó�Xe���&Weo�B�2FC&�:����7w�\�\z�g`��nY�;�la����f��-�Y��GTep��q�u���Ӡ	F��:�:15Q��R@�R���U���X|E��na���5CH3����<h[ǥ	�}�0�JP�vM�`��)q[Z�|���ۿz#!�1IaSq��6��m���c/i�����Y���Q�%�Nb]�(��$��"�2цx<�o�܄������<[��4��h@�ǍA�䋊]�27�M��kl%K\2����9���s�d̤Ar��h���\V1�O���K�	vF������[O���I{��p��W���0cV-	u��r�`%�u����4"4���Q[J�}בofb���oS'��ղ��� �9N��oZl]��$�7a91^<�p.R�G
�-B~���}�Qe)�sj��8�_��j0zCүԅO{�7�~�yo�Ԫ]qF��7��~BӞ0��	���x�5ߛX�\���O�C�U����Dh������@��W���(��)��J����AR�9Ӆ%%J�3؜WL2�Pv��X��"Re��4;AJ�J)�����I���ͥM�� 1N���L�3��i3�"�7�B��Y�.Œ�q�L��|Z�M<���9Mm��%(Z�W���t�Zh��Q�$v�D(?.��S�����z����uR+ެ���~ua����Pb�0��Q��NXZ�����c�qy�{7�1w�4�,���wt�3��6k��ˇ�����#K�D6ܔFeu 
n��f"�*R+=(�J�MfeP�%�kl��vw;��?��C����A�#�[/���3�Bh:g��Ydī$�Ƞ===�y��V����w#kKN<���ս��Й�|>,��gI�2��"����o�+�t��9�^��S]���[��0R�pŦ�t��w��*���n�4�&S��!��:i.�\��ޖLyV��x�ing:��O�^Xl�����.w�X�ꠘL� � %�>�dӨ�T&=� <���k:k.A3��X`�������mI} �����M���o�rW�4q���l"�����+�Q�MB���Tq�D�R���嵓|ry/\W����B���t����ۨ����ڕ�cOt�w�#��s4�H�5x� +��S�{�@/A^8ddDE���³�UU1�'h�{��pɢ��ǫ�%^������t�zS��L�j���6�0�3k���z�������\n`pX����3�B� �8���B�:_A� [�����S������ゴ�w 9�L���JI/��eN'���O�d+�k�~��{\lQ@J�ҙ��ɚ��\����or� T��k�h���B���]y��@!����cLB[��3F��1K�l���Z��:�P�7~2_��8L��c�A۳`�aI�d�x���\�)�}��ߎ0Y���s��+5@ї��2��v&l6�� #=_|�:�R���@���XD��BȐHh�+�45�U��b�!C��|�s.aQ[@�j�Rp�VEi�����}�D�����,��q�9;�Q!V�>���U�#%����s�;A����<5�%�����=y/�SH޾�Ul~E|���R*e|�ˍ�Ҟ1	n��܋b�@�H_���.�X���1U8��Ƽ1�%E���r��i��U	�A�Z�V���w"A���ʰ9g�h����勒��D-/l�'Gaf��wM��B_���r`FY�e��Y@�����;C�gn��͜Tuj}<�F¿��s��dЛi�Tc
�)D\�B����l������>p +���u_�XG����碌���#���j4]��"��Y�qBo�����H��&�m*���f��?��h���9G�j%R�#��2Q�#�<L�\"��/��g��q��D�!���hڜ���u?�� �'3t9��]�ܗ��&x�KP�oJ���l̕�L�>�ɴ��^���
���.�������k{n�Bj����og�*|��cK��ϸ(��.����pO��៱q�^~^��r �^�F��!���l�Mx<�I�"�6�F�11�wn�Q���c7�A}��v�TM��Z_x�
�:J߅%f��i��Xν�C�N��x���!oꙣ�-&<�/]/vIN C_6�C�]���S�KT-�(ʓ ��#ND(�#�d�������`}C򦪼����^nz��SSy�V���#�|�^��!3�§�M]��� V7��ڙ����2ݜP�z���r���ՙ�3���)ٺ��R�Kp�u��4�r �Lt��^U �+Ml�G��h�g�bL���Wd0�D
&�PtxѺ�e��L#]�H�!�o^��[]ڿ�Jd"`�#iPu��lU�Lmj\�QB��a*�1 a��z��w��� �(1q`���up���uR2��K��|�t5��eG|J�oAj��� z6E,7��QA�)���)e��w@��/,y�]�ϣ�5x��}6_�ᮇHWP���c���ac�Ow-� s6�f2�%1{�̽)�,��=|ԙ��\�E'���&�Бii��guP�F���Rر��a��n�7�p��q����R��\\I��]l]�U��V�m&;�
��$Av��g��^��*6��'p�;����HX�|
7�g�P�^/�8�g�%�1A!�& 	�ɨ����UN$P+0�8�}0�L]��݄s�3L��&�me�o��O��5�O�F��t'��h	�^�k�q.b�Zd�����5_ɲ�D����6.��p(6nS�d
00������Z�Z��2����2�}�BG2�-/��3�w����8��ewĶ�11�JTC��c�޶c��	��M��g4����Oϴ�%��^���"��x�/����_PK8���d��A^=(%��G����>_���?D�J�t��6�T���[w��y�֙�M[�]ݢ�ED�\�k(�QA�;���oܚQ!Y�c2s䈓i�4���}��Ѕ����$g��*�(����I�Ɖv�w��g��SM�F���򂖸�
�N�/������f�3zF���xCa�p��u��KϘ��Jh'�v�+��^�/��R�!����ҠY_3���A1����jwe.I�W|:�G.M�����+��cdN<]<eE�e)>��\ѹ0� ���0�S���t5�㥠о��$5�ӈ����j�J{�H�y��}�qjx��n%Ju�o�F	��=�j��S	�Yj�0%F"+�~���	r���E;0 E��9�9�H�\t@a;Kev�h�E�<W&ڮ4��(oE|g|e�dD��'��e�d�����#fO�`
���Y�/�"�+bBW�"�<Pm�V����HB!lF�{Q�C?���RW�L,��n�?%�!�|ƌ}ȵ��U�6�J3i�`$����QO SQv��Tl}q����Ev�.������a'�큊a����K��t&va�؊S���ӭd��<A6�z�	�\�8�c��wH#7�RORQ���ٔд���l)�Gz���Κ�
(;�@�j������/O�������C�Њ�>�>��&PW�0�@���O��P�4*|�0*��>�Y*��d:���"{�@����}��� ��0U9��9����$��P���l�=g�>} ��nS�ǋ��M�� ��6v�~,r5��XZ�7��-�dp�d��\�b�d %�%n��`;H�cI�B����3![�Ȼ�T[�[��*�|��3"3 �G/��QO'�iڨSZw6s�����M�j;�Rbg#��
<v;�m���v��0C��I�iο9%����ns�)����n'�e�ݷ�ʥ��lR�$<:�f4�-4̮�N�j��J�x$�$F�����?٥b���Kc��f�UF��*ЁFQn�a6.�Q�he�(ڸɇs�6��r�&�s��YdH�8#f�S�}�8�^�|n��5�_>td�{�Rб�W���d� 6����+VI�/�c�5D�ޤĳ�e��yu� ��<Q�g[y����HzZD�W-'9ɕ	[@��[��
�\�z3���!�ތӗ,�9z hA�'YQ��t�{I�-<NdS6����$� a땮�)�7��R�-�Q��y��@B���|$�����r��Tb��ܿ󥶗9����t��1�_���裸�4S@d�xz�x��5X��,�٤B�XS��<����AU��{�aքU�쥨�x^=i��T~�����y���,�wL���#D�U�iB�\��d�%�<���TїB=cW���F�d�Sf%��g�^#sǅ{	�Y/�%r����{�O�,�� ^�W�<'��J��}��G�x�{�Hn��D]��?`�Q����;�U�Q>��kw��f>������ɰݐ�IYó52����|xv/�9=��9�����1{vDz���c"��Q޻�7�t4�<=t���t1�S�,~pA3D2i�s?�K��������p<8��4�Nt,0nP�G҂�1��q���\a�r)c�Iz���z�tZ��ys��[;�d��(�\h38�-斝�st�.0~������muZj�묪��]B{�3�ߎTM����pO�����U�m?�� 9hh��N6r������S�	��T�����4�+Rv��O
��9}�͇���  ��E�r�{g�
0H���T`�./�1-��6����<�*:��x�|9��o����ӒFF(�[;ＺP ��|@���g�F�#����z����J\G DL#�f�ꓮ�;��1Y+�����g�~� >a��l)�E l����*��WV�|#��H}o�Q^şJ9M�`J�- �5ʜ�I�����βY���7rճ�Ɩ6C[�>��2��<�DY���"�g�#|xօ&P���ܥ���9&G�>Iz�
2���6�@�� c�3�7T?�a�wx�mz4D���@́Z�"�δ�$� K�>��k54����jy��zm��I��$V�Han�.�9�� `���ɩ&,o6�}��)srې9��46���P
�]�3ҽ�{j,�0�`���+}�ͩ�<o�E��TS0e���ߕV��,�D�V�@C�����tE��?9�8`�kV�@&_�ʫI�){�D�ݎk�(~��ʓK捓:��K�4�����G�� �,�� �`����T�&������_eX�N������P�c�<)��?�
k���0A��ɥ��H�p��p�7�QXV'�L"�ټ�.���a��� �f�m�0�&�0�>k:y�v�[�HI�p�"�X4���f�Ϥ�c�R
o�m�YL;���T�hB�����V����n�� ̮+H�s�m��g8�y��:��8��th�Z�1.���t�*�p�/�5�%u���|��F�j�=[Pd��1>�W�d�!��1e+��F�>L�$�w���4��@$�W: 4��P���[�$��A��D���\��e���^>�������Z��_4P�wɡB��@q��3B6�.����)H�Uv��{��0NaC4Oc�}��f��D]7�0�M1��O�`��kx�X����2?$aI�g���`��`���|S����O�N���58<$�ۿ�q�x��X
���2_�Q�K�t�>ګfOY�**A<�0j�c�˜�h�S��D(C�)3��T}	����H2f�c�r�w�s��lɥ/�]@	i��������&˯��J�i��1>T����rH����Q�M�d-N�`2����5�L���Ϳu�cx�%�i�-ѸǦ�c^[���Z���Kh�z��@�����J�I�6��;;;�<��E���iH'�?��|���l!2�0V���(m�[����b�ʅ+�+��	Ȋ~Nہ��d�jc�)xb�-����|��U��ej����@vb0%J�/[������M�^�2�d��Z���,�Pm �`��n� p<�ȴ�{�̜T&3�ѿ�8<��s���[W?��&~���h���1g��UMؖM��\�x��c��7��Ŧ�Q}@=A�K3:��#0��V��!>�t����]
Jq��+>�ZPZ�JḤ!�)b!�`C��9X��^��+j�4�F̨+=*$�!!X� ���A~�j�Ո��_"�}��"4�,�$�[����]5�1+��O��] b�u=r�(J
�����֣�h��$�HP5�,\4�յg5��`�*�H\�����/^�+(�.�=;ۓ#خt��xSA�U(u��5v$a.� Sqt���L�Ws�u�2���6��)���/u�U�K�j ,К4kt~~�L�RJ��V�cg��4�Ei��,��Rf�gt�I�%�^
kSݪ��Ay~m��)��YQ��~�����i�1F��8=Z?�I}�}�"���(��İ��x��rg�G�F�mT^:&=��o!E��'�b�����y4�+�g	\1�bM|x��G�����#.|]����hJ�?���	�����h��H/�T���
5���1�8���ٔ������WX��vs��8^-�oz-���DS����Kc�G��Pjo���&�b���*"5�! �L�����t�qPe5q�y�|��@6�����Y,P1�Rj��h�J�
;"�����n#9����eN���*%��#���K�D�<��TTۋKl��8��T�I�M =�N&M������'������|�
��<���%=�s�R2�H��A~ '{Í���4F���g
9���g�A��?vFq�t!���IN��I����>�"H��`zC#�O�����/��ܖ`�]>��0�9��9"&�h���1�3_�+��R���\\
�K-�=���<eɥ�e�U�SyZHy��N��$I�w�w��jJ-B����-m�d�|7-����G��#I�х�N���&d��I�²7�ln����'Z�����)75�	���	H#�R \�ۤ��ش�D_$�'��~��*wL�/<a�1�����k
/�ք	���v�[��q��
����s:`N;�`Λ[ap�)pӲ�����czH��hl	�^�H�b^�IJ(`��n6ܤ�)H�C`�ϣj�:�<�dMP۝W�:V!HC�aN���/�la,�4*�.R��O��XD[^��ߌJwx�&f#�a�į��{1�X%��S�B��/#��.x���g����E�-M�F�_Ah�8©��O�$�q��BÐ2�4E�C�Ÿ�@�*�?v8\��S�\`!�3vmL������ 0 e.��1[�����9��b;�n��!����hy�d�R��U�&M�I`,ZH>T �]���'��`*����U�ϫ�xƁ�x��������3��ڽ9s1u�����0��Q.��"nL:O�.�/�-���tb���?����	��Yɐ���6�wT�v�vE�x�F|�����C��CHXU� ��UP	��6�~AB�QȥJ���y��8��qzB����F�2�G��@=�L��y�k��ORy�ԿA�t�R��d$�_���.�ײӘ+a��/J���w�y�3/��\Q�Uީ��B�,�������� f!�LE��&��}c�Wh삞��V�Z�\(D����t�)V�V%8�_������~(��FB?�%������~ƮnΘ����oi5G��iM�etc!�a�ߋ+?Onw�s J�r�"H�gnx��L2P$�f��r��h��cl��Շ��ĉ����j�EN��{����∫}
?�o�TS�h�@�kʞ�wJ�~�O�] `�0���Of�ҽ����E��k��;-`������~��.��"CM`n�5ds�0;����I��=��;1k��p�H�k��O�
H��B����{d�?0o�2�\p�����n�b�R�_+�w�ge�Sv�*`� ۭH*6�q1�	���rx~Pq��vY%�J+��Ҧ��`'�Wh/���G��U�4�^�5I���˃(80����}�>9��$�|*�f�hτv/�R��PǠ���Љ2��}�,�],k�L[|���\n.0��4�p�}���8�������Y.�;�p�|�0-�~�}.��y�P�h�e_(�󪿚g�3$<b`�B���>P
��I)��|�����:%&-DV�{X9�9��7�k(SU�9�Y��Z����m�EKP�xZ�.�;OZ�5?��Ą�c�:��<���Ժ$��9�0V򢴇�/�� ��c��@+'��!��N��m0d�/)9�R)P�ąű���I�?AQ�!���-�
���T짲�ȹ��gU2h[�����:^�{�7�F��&kU�߃".�<��[1�W+�X]��]�<�(��z��x�����h�P"g�C3QU������a��ށ���w�L!/�b.��V����\������>_!gM|Z�1`�*R���RM��[)���r1�'��5�L�wǈ��:aEG[.!<�!hK�<���U;�/��5����S�m�F�G��7��R�r�Hh���6�SŞו��A5ath��]�K�:w�gص=��l�H3��-[����)y:�����!w9۞"-aC��a��f<9v�H�{��xU�.���GF�,�!�ӥ���y���F=uS���N���e�$*�݁G�܁�2��e���YGQۦ�x��B���<5��,t{s4���:%�ԟ���c�*��{l�8�����Y{�4F���g�*�,��ӽyR�y�F|��^������E ��Kؽ�)Ov���n��ܳ�N���Q:���b(�n�ϵv�����I�^��������1�#8$�?��3U5���S�^u�.���T;��1�⌖����b��G�)5��x��3!�x�=��=�,��C6)]n��p �	�3���Rx�lfe�4���ǟ�tr�e�@q���f!<x�/ I�;m�a�b
�A�?�SZ��9`��!�l�]�dn�+����.���� �o��ݰ��yr'C>��j�J�n�צ�&�#�ls���$Y*���c��
��Z�x�Ϋï����E��N�z,�)s���jly%����1�����׈�M��pg8r�+�Q�~�BK�|�h�T���[;�u�-&��vD}���/ �.vII���U��#P��N��t94̀I�F�Rj7�׹پ�g�����&G�!!і��U�=b�:���\)�cK�4Pʐ�8[ƙ��M�-}�J�uS�<磱eq�=|�����l�b�j<���[3�_9X�ɑ�g��5&�'�'�F��c�`�چX�v��1�]�R����ژ��U#9tj�M���[	B3ȿޘ��K�x|��!���겿�	hׁԻ.�]N�C��W/�⧃��F�+�Z��2D7��$@`����呣�E��Ĺ�|
�c�>�kE�f�Ŏ��EG�?eN��`ǜ�
5�@��ƞ���9�]*k�Ѵ𴶪�\��,:�9u���|��'���
6�E��K�х;�=2X�\{%v���a�T��;���?[os�,4��$9�0;/.�ݚo�(Gy���������/��i���um2E�E�5,c�r߃���p�����#>�n}ַ�5;ۄ���^����>���Alt�-PY?�I3��MՔ�5��s�;�����\Q}�/:�v�B�(�Z�ig�&V��>��o*~^(*�o4��×��	�hCy֎��4��w BtnX0��h�fQg1��`���[��b*�H�A9J��'C�_\�&=R���"�%̉�A\�i�B����<��m���#��q5�����bP� �g��-,������� �H 
Vy_��kBLb�4�q��\r,�J��kw�D� A~oD���KGh�q�UCt�`��2����'�'�8ߎ�G/*��O6L2J�����΃���W�L�d���>�u�z����z4��/�g���Si�@��tq����K}�������.�&�̾Lw쩂 �:���Z��&5G�Pr���	
*�9���q�F�A^��,%H�/��k��~S@�~*�<��6$x�)��b���!����V`��aq���\�E�@�o��j���9mQH�w]z3��ۼJ�l�����ƨC�_��I������ё��W����S�M<�А<9�>�U�P�����ت�M����>�ۜh ��\�%k^Jޫ�٭?7��~oBd7�a��-<&#�2<�ٙ������a=z'��?g��^
�2˒��L~F2�����Y�����ڔ=X5�~F~{�I�XƘ�8i�*�gR�7Q�L沈���r��2���}���I��7��,cm\)���|���PK�����hlF=�)�0�xs#�oJ��TҬ��Vz[m�{�as/�s(��c��D\<�׀1\����\�p����3��_�(������Cߝ�0e��� �@����n����O��>�^�{gz�~��]�Fx0�>L��7�v��P7��s�ǰ����AZ��V�3��Q�)ʋTcxѬ��~i�N��}�Y�Á�C��TO���	�VÕ�]��g"XL� ��;s4D��:�>t��'&(:xe��������;��tW���>�캸�t]F��CF�T����_M����l6m?��� �2�^�}3����(v�8�#�/���Y�tYז<��)����5+V��~.���ݲOL3�q]�Hv�P��q�� ��]���HҶ�.���pg)�6�3f���1�V@
k2(��i���+P�Nc����?³�N�����Iz�-��ē���jOQ��z�&x��(8%����#߁�������"K`�U���O��ؐYfծ6GphsD�$���ݙ���œaG�����0pd���J; ��A+��nj�5q�?���s���l��@�L|�6N���x��|Bܵϋ9����8}ė#>�� �F76Z����ԁ�t��{l(Kx�Y���67�jN��7�|��72I5�Ie'������<��={n��|v:�\� ǨO��r�����6�k<�ubZf��EՋgT�}9	���V�L�kM��'u$���Y�e�
�>�=����06�@�}�O`.�Ǫhѽ�� ��n���3�@e8:`���If�[��\���"��x�#[d�0bY��A�6Ԗ����������
0�in���m4�փ�OթE��4���l�?+U�
]���5��$���$�Q�cQ�ʠq�/D����GK�Ј0�	���Y�6gy�~ H4��@�7+��IٰV�U�%�S
yq���������g`+���軞0��=I��{��Yp�3M��	�]��M��8C���'���X���hEp�Du��kg|iW{e���G���΢�.zLT��~C�]] �NV��)��R�P������@o>�\��P?��'�-V'U��,�_Y �O��u]ӣ�����?6��Ԕ/O��䆼�)�\�k���৘n&��F��VK��(����c��Ҹ��T�?�1=cq	,Y?�8���Y���"0�����+��ܙ�㠧0Y,�E`[��'n�Ѕz����5P�ᤣTfRT��{Ԧ"�K��z~����kz.7�(�A&6��P�M���٫�"�m�S�c���OP�z�M;�H�u��}�^��,-���RU��`u�A�-�N����?G�--�k����ǝ�*a��~o��&e��M/N;���g5a��;��G�6����9�%����֥����:�e`��:Q#��y���/"����(ļ�2�[x����Ÿd���I�0%�֊T�P�#{䙿M"u�u�JZz�`�������\��H�r<?���:�[�T�|G�76��� ���oG���L�[�CnɁg8�t���
���_�s�����I�IF�1��RH�6F��)y��_�R����W�m�|,:�7���|�׌D��\ä�CIX)�=�l}Hz�l�tn+H�|})+��O1�CO��˰5// �����"�:��w#E��y���l\>���
=щ^��݋k��9��'����XB~��d\a"fa�	fC�ۥ�|�?�m��iR��C��0�X.9�����V���`q���0��M�x��=/i��_�,�dh�w:��O��@��t�Ba>V�.~1G��A��pbI�
�LHl����3:Sw�h��|��7@_��J�H��{������/L���X�5|���k���?$�e�80U4��/�i�U��qX�%��(�0�R�%��7b��Ǜ�:��Ц|;%JtG��`���<Mwf�ݛ�VYQK.Wz['˧˔�=��ەfQh��P-�k/��R�Sb_9�8����nVDc	�Ag��T���S_��LjIx�A�8X/��;��u؞�2l~���5M ���H����Ov�%{���ɪ2�E\8a|���Q�7�f�4�c�W<	5�D�r�_c��8n��fRd�?�q��"��������*�E��Y�Km.�v�^�-��_�!��Өz9#L9��HP����䰆��zEѲ�����#y�
��%*�fO�+KT�������'	tox��<���dq£fI#El�YS����Ht�տ1�^�����7�)|W���-�ފZ� gX����Eoc2=\{~7�Ȗlu�$,n�)햗��Z;˽A)�X�J����]4��B<��eD��mN6�^�%{L_�t��і���i��^<�Y[S�����ۺ�Vֳ*E{T�F *����⩲F
(�ov>h�S�<���-Olfx̴^?�ҋ���西�?ˀ"��0=@ �pM*�<�� A�ց��ҍ��"JH�G4�5�c��6E���]�Yo���mD oG'J\��c_�dYFao2��bB!�]�|w=ז�X[T0���� �Q��O�<<���_| ���6��O��e�;�~�e�f咂�Z���I���Cn/�-&	;��>O���� 3%f��D�~4����r	�H���T=�rjP�40���x3;y�NJւ{���V�����Sڵ=e��5��C�ߌ����(��&�c��GXxm+r?�~�����2�)�=�[r�(D+b�ejr�����+�#+�?Pǐ����yL�U'����p�2��T�,�<��%�eGa8�O��,r��*�fb)��$A\�޴��{������8o-6��g���'i�vj�@��Ui�S�90}�{,T���pͥM)~�qµ<�X�9��Gvgs�R�*;1�CnV&8�R�Raaꏋ��Q״W�g��,��K#��M��̲�R�<Xn:��Gy��_���d�y�u�����ehĂ����R��\;��bW�Ѹa�71���ޫ�Mahj�)���q���sg�v&*�Q���e� �p���/�@���*�R���$/<��5�_��{�,���ξ*�B=�Q�h!����$����9��R�H����J�>�T9kF����zצQ�*���4��|{*�&�4���I�;��m�P�k�U���%R�����6��:D��B�J������V�Ӻb�x]+�1X���%mm�D, _�t�FT��bg���v��򝻺�q�J�'�'J�V+"��[��v�܇�研���c�v�|}�ﾶ��$�HF�݅��Ӝ�������T䠢�rO��	�&���#�ݱ%5T������~��� �6��g�� ��c����XMfa�ñ�� �	�A,��b�%���$��D�9��2>g� q�N�`�O:��?�{	H�Wi=:�4���An %,��V ��
7��������(a����e;�� ��>
�'��u��T'r�a��1�}��K�]A��N��juU0Dg ?B>^ܝ���U�+I.1|�9�+e�=�=!ߐM1Q���fV���f�>x4�|Z�}P4���D�u u�K�h�E��sk�
�}^�Eq<�̰:ŊN��E<��h䮖�L��"74�w2�v�0�:T�1ӥ �������;�~���`��ߌ)��@�'of<R_%yv� �$e�*u����C��3��J�e>��`������T�,���s�$SO(kd�Fk�~;�A$�O��Өk��n~`�sJ�!�$n�;m���ɚ'MF����V�UH_<y�w68�ߠ;i�Sf�g�8/I����6 �@�yD��B�=SYL�kֶ��I�D0�"�u������=�ep��ٻ	�i��e[��8"���2�z��12}�Ӱfh�00�|3�=!�����`j�$�����k<f���v�9ڂ-ؑ���l�H���s(�x|,>���Z�S�t=�<�.��uX"�D[!ޠeY��M�D>%ᦦ��������8���T���7�Z�lĳ����{x�R��I��<��m�	X�Iέމ$������%Hƾ �4�
 �(^Y����������ThGIY%L�u�y��|� �^��:^�����n.ǳ�Ε� �0}獷���rX�����Ub�P֏6q5%k����W�W*���/�/{�#S�%OOu&��� a�L��RfC2P�������:�4"0�W@t�ew���֨����W�3��ԙ��|"��d���튬����x��9���B��nۺ|�V]���� ���3�a���K�&儆ie�HMGN ���Ei�`���S%2'bD�f�k_���e�'*�J���0{R����SX�nE� �"���Z��?:eN헄��)�wb�"���ҏ�?��J��M4��;��zv���N�WH�{���{Em�*�Ø��@�.|�3�r:��Qos�=�9p�|J�y�oGw�t��B'��J��3�JB��&wr_٨}��z���"hq�8�� \Os���ʥ�DEy*�>/B�.A�~bY��u,7*�
_'����W���5pF�j#Y�s�):OEv�#��}� ��K� ?9&4%��/�U���Q~�_�����r���	Z�Z*U{�F�Gde��N����q����T����/ɔ0 o�@�����r�/��+���0ڒ��*>a=5[���&��޻�qf��rCl`c�#` A�k�5��w����AP������`�������5�*&IJߓ�Q����7�
��&�a|�	T�qK����:aV(I}�7��Ty)�!)��n�H��rr>�`������~�L�+k^���S����
n�J���r����Q=~h)(�Ȭ"��+�~]�F���B3�\�.8w�\;�Psf���pη�N����(mi:6��)�9��f�z!�k�-�%��0r�N���^�/�!�@���z�	Mg��x�!/�.�
. ��/�Ў;�(̖y%�q��2��ڢ��`-�O�����Ǧ,��X�.
p�6�ah"��7`�(8L�[/�kI#�����g���Ϙ�(u���r��93�w�<��-�e���6��/>���;�sˉ�{G7��~BM}�������Go�9�V���1 ���ќ�N=�o�:S*��QΑ����$A�D�T�-�S0x��:>F���Y���TloM]E!x�Оz��L�.�w�e���c��˽�jA1��ː=��'o���1�5/rMg�I����ڡJ�`lH3M�.�4�?�|O˔�P��]j���8����0��<E	�Yz����_5��W*��Cq*��@�4õc �Z���u5�^��"�X�Z�s��T&��E�dn�Bs�q
T�İ�Mޮ5�?{�R���3�Fb��]5��o�S�Y8؀_��`�
�C� ��8�ħ�BX�Ũ	���B���wgѵ׾�B=�q��6f��H�̥��f�(�Â�b�z����]��A��"�\��;�GmzC��?a#Ы$o垣]ɯ�g]q�M�#��$E)�"d���y"�L^���Y߷��j�%���xr��4�lm1e	��ș�F��F]f�c]����i��s��KK��/4�\���Px���i�J�qX�˕��zMt�X�%�
�I��xj!��~�Y��:��b��������➣�R٤n(�|H�Ǩ���L���C.��:1���c':�\�nl6���@�٭6-�J��뺖��`jcǖ��]v�g�7W,�k1��~˴9�]�э��ݢ�pW�l�^s���V����v-��c�x������=��䚪K��i���;E�wq8V�U�OD}��wP�������%��Y7�1��9o�D�Ƚ$�.�-y]���`i4"s�*M9F���ܷ��XE��`ꓫ`R��@���d3ƹ�	��("د�����>�x�0`�7��� �OF��F���|̠��Wժ�K�a2r�m6��_���o Z֟D C��H��ck�	,@Yi�O����FY���.,�;���j��w�%|��(��F�mTV Z`m�(�[�T�vE��|S�)�X����q����>A���#$U �׼Ki��H �m��H�\�����l��7,)��qۗOYY�X7���ېܶ�g�k��j偳��ƫMEV�&<�Z��)N.QI�X��5M
}�a�Ho�|#�)N���L������I��@_p���V)�m�i�4��k�±�2
�~{M���j�7qt笚d�;.�"%��f�q=�s��ʆ��i;�y�LF.ջ�*��%\�{�uCajܽ;��)�}vvS"#�}���x�,eJ덋���N6ܩ�`�WAy�y��լ��w#|�2[���~ �&h2�o�6��+ �(�T�J���h��Ek���a�@Y�H���^-I�iG9]�TC�,���|�XZ�/ዲʋ�T���8�掟�w%'c�L����0CЯJ3L�M��X�b�V
k��X%l�ϙQ�S����e��}<��W/�O��P$��a��R�ͮ_�h�
��;W�X�BZ= �����5\�ih*V�&��� ����æ��ǧ�&��0��C���4��kFgI�?�s�|��@�r������#��פxjz��G�t����:�o�in�*ο`_n��P(TDq�t�!�;V����:]h�I�)u���(U�����N��D��mE�i�e>�wbQ���b5}������3h��M���G��k�E�~/�(�Η�e\/b��Á�Ag�%u��*�kb� F����yf���7�r�#�H��)�⒓z�ش�1RnF��h���F!����P�.����5�T�������2CKի�k�m���bRL���y8J^��_���נ���6�sPΘj�s���C˛	X,D��k��si�;ܑg��+d�����Є��>�� Q	ecb�g���}z���:S�57���/F(*=4�L��X,���B)�IjN�����$T���	J�K��|��tvs7�nY�#�G(�͜m �N�e�p�N�������#	��U�A˂�`[:"��&�3sFh���Z&�S�)�����~�3�<�?aHDd��?[�d
(\1Up6��w��p��Q�0�b���A���P���NVHi���v�C.^fi@˖RX�{�s]�c֥�rM���c��	`���#��~'�Sh��[@��bU^A Ǣ+g,��Z�ּL��UXxIH��
My+�^����qƆ̰K��܂������^0��>�Ƒ��}���u}$�h8OWy���6b�c\��Q�-�ݢա!�l�\j�f7�����P~J����%,q�㔾�z��'�2˧q��i[e���8r~8��C�����杴HR�I��Su^�,��%�	������Y
H�̉=Z��__)�T�{�ǬڍݼgUY9����L�W��<HBb𲷷���2�7a[�*y~�֖+C�X����o&�҇,lRƀј 	�p�����?��c�l�~ٙ�0A��(���^a��r0��Ն?��y�UD�'���_#ufj'�(��NZ�z%S��K�-�û>%ز��z��h��<���A?����Yq��xgUa�:+¤A�5gDc7��/�I/�X��J��o�@�Ld����8�O��9�9c6�-u���Q�H�a�� ��F�`�P, ��82!�v~�G���!"�
���ڵٕȔO�?��q��,��sU�2��O�	�|mk/+y[�uN0pji�j���}G�^>���2ݸq�a�t�V:a񢾾���)�j�\�����W@&
bt�Oݠ2)�{5Xݧ�Ӹ���C��C�v���W��v�2�"����S�i�es|I�{��K���	�h���hr���t��!�zH��0=�錗ū��@�L�6RK�P��1�j��ao
��L�Ƥ]ꫢ�V��a���*�cT�i8KD�I[f��nk뿸[A�?��(4����m���L��$5&��(��r��L�y��AՂ�!TL�4IK�@6G������~8�aT�U�'���]���H�=�*~7%mtX�����^P�mм7N_î��S���h�0�0q7�6�v����a�v���86E[K+ۑ�������n�Ͷ=�{>�0D��J����Y��U���'�+T\��t�)f�����l�=��U='��n������}샧)��4�c��Q�jӠ�Nm�����XBƮ�sV9ud�W�	Q�����5�Ț�|D6FU�:ap"hhhhB�G�gE=
{W��/��Ҹ�Bx�^���;�is9�m���%�:'�Ѥz�'4�1N.��H�F(�� ���ݡ�����s�B��QX�_#��Ё������C�٬y�u8ݒǔ���[����}�[-�v��v��Eؗ��sC�w��pO��O��[Ee �[�$
f{�>#1'���Yņ:{Gv<�nP1O��f��5����q�I�Lb�U��J0m7����`㺗�@�飄n�39���BF�:#�wU)����oҙ���K��3"%bxc#+z�oY�~�+�/�+l5pB֭Y�0Pm�-`S��w����	�_�0X%7ˤW6�-k���Q�a^R� �%�<��9x���r��Ѥ�l��j
��^C�����Pl2�{WA�+��RR鱅��fӓ���T�� �aS�k�V�ѓ/�7����=�XHD'�+�9*t�]�����;��W)�� ���_�6�z�,`ms >�X���rljv�aT�����������f#�l�}�"D���ƞk?PT
��C&�-�A}`��ƕـ�1p�7 ��Ѩƅ��+H�x�p���h���gz�nc����(ق5>I���ME�����Ot;CŦ�F��5��$�4��U�1��_y,Yֻ�p�S�'�hq�1��p�# d��Lϑ��+~�W��c!g��!�X\L\IXE����N)�X�L�l= ���G�N6�-�Z��eT%�@��3���o�C�@'ojs�����s���./Ա�S�g���䯹i�5p�5�ar׮���Ϩ0i2$�J��>����V��cq��~\^��/u��ـ�u���u�^��1e���u��%r�34�[���|�o`�aU���`��^��ǽ��֮���<�U���ws٫�d��h-O�|23��c�u+$��\���aل����Dy�k��@۟R�Lk�8�Ǘ����g���CUF��k�l}��C��R]�2ŝ�8��Dd�l�������R���l>��=���/ J^w��4���!����؈Ɉ9�|�wR�[ Y�6x6&r�����D��>�Ԝ����i�I�&����Z�\���+X6����Mu��G}4W>q�3��>�)z����l?[��6�)4Z�h���y�K�����ƒ��1��݁kNS���W{�f�)��>-I��@��Z\��h�2�|V�{��=���AZ�g  �D���:e޴�{�c��@�!��KZ�v"��jf�2D�������F���~qG���$za�p*���*b�_*^�]Pu�F�=���j�a��_$�kA4 U���a1M�J�d~&�q���Oa�E@�Β��K��L�gAx��Ӈri^MMp�kQZ~�;�Ni|2jǕUu�?o���J���k���fӀ�Տ�0� j�+�Ye��EE**�Q����_��t���6{Ᏸ��z7nW���v��>��(%4�|:#B9K>�{���5��0���f��čz�3g��x��0�4f�\��`̡��ҥ*�(��U�g�-.LWem�!�!� ��$R����)U����7ȵK�S���C�Y�1��WA���@�;D3�E�bq�W��]�θ7r�a8�)�D�F%k|�Q������������Xj>���"�q��hD<O4e��>�_J2����t����`�)��%[8}��E!�O��>qh�Sީ��m�>�9N�݉k΢���4���q�#]�Ʀ�\�df�@��*r�U8��h�#�Ķ�Yx��^���H%��\7�@���4ђ
,q��_/�%+]�6��|��:U�`����T��@"I�Wr�Ǐ/�*fʫSu�y�����T�ކ�r�f���R��Ę�.��{'�
U��0m��*��5��k}>�C��	�?��U��~ ��?�{���d4�G��DQ�2> Y��e�.$5�ԭ��ěg�Z�3+�2I^�0{Пű�G	dD$���j-��y�Y�X�^
��n�m��aU�������2��<
!�2�U���6����Кq��,�H�U}Q:���n�}������\q>t˧�Q����w�oX�yJƮ�4y�I���y��$�ܿ�>K7QN���-��+��x7�X�U�0�+�n㿯�ۛe�q�K�����'�*�����QO����t��lz`�m&��#z�����+@*杣���쬮ܱ��~�MM�?��[�$��|j��	�h)͹��vC��IJ���fCg�߿��iT
�s���<KO�xK��C�(qCu�~Jb�m�����i�1-R���c&A��W���AA'<1_�m�Y�g��/,t/�1�e�=�8�y9�9c���}��z�fͿ����=R8���~���4��qI�����e~�>���]p�Frv���5�3�>[�i9�}��T5e�F�)Q�~�hmy�*����������hA��f �)	lvZ�)?�T������B�,�ϩ�g*�p3x>�4����[L��w�:"��;�1/����� �GZ�s��S�����`Jij�`��� /(�r�_��S��T�)-a���dW*]��\��C�q7�ki�\LP\ �ng����y��=�b����`�ǵ�H��
WR�#;��O���ķ�&�ک"�vx\��H�6�r��]�۔��v�M���$z��(_jwwX���@��V�R�q��|�_V�m� *h+i���1��0�4����;Z"�䋸9Ѡ\d�hm���d!b'GV��C�´ۖcf�-C�����|R�J��<L���e�vU���9��Y��趙�iG�!��Vj�p8p��O£�B�
##=��v��)(�־v�_+V'	�h����Q�iC��3I�&���Q
��)�?��8M7`Z�o$iϙ��bBx@;���5_ϝ�U�5M(|�|��NFNZ8'Y�s����jP�5v�|�-	�ͷn)�5q��,�3�#1����]^�ϙ"N]e��G��m�.E-{�m�4��"+d��9̝{ғ �wp):ʥ�04��ܤ��+�_���߇ςI�"���r�ƸF��q,-��8��z���CwYA<��,Ig�K�|��w*��