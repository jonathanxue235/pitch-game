��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C���7j���Eb�Q��gQ� Q ��������˻X�"��ű��\t���@���痄[w�l��>�\�_�w�W����K,��r;���Q<#([ۂqRs�_��7+��b%�(D�PUL�++�(��Ow�Ö"��A��!��]��\�q�t���y��]�ȾuT����)�;��g�*�b�GL��X$ʾV%-k��k����)��W��+�a���$N�EY��kx�o��B߳Q0��|�(~M{�1y/ ����'2\ː�s�*Ӓp������iĺ-5<֌�I\ť�U���G�v�������Y���Zѿ"�kb<W&!�=W�^�*��';��=-yk�7���Z���e$���aF�I�(�����Q��q� /䝵d=��	L<&"���UN'�WU���u�
�@,82O�cJUs����	$�heA�Q�����&�П���	_i�9�C����
��r���3�ug�R�VD~r��G�5aZ�ˋ���a�����l�ޥ�Fr�h��0i%(���Tw/ �^o�n*p��fq@�Y��+�+���}��ŝ9H�n�r*�F����c��C��SL����h6��4��>��[��c�~
4
4���JW�,��B&�������g(Z��o��yV���oҬ�5m�/� u��M�����8�j���1N�p\i	��"*Td;��s��;"hE�1u�,a�.p7�[�� D�ށ�럊�[�
���2���we{>f4�-|܁v%3��M^�w�]nj���>����F���o58�1g�4��%�V��%��a���G����v��M,*?o6����:"u�+]���f'����Yߢ^ь.�w��6�����!4�J��eA�o+�Cj��}Bi�r�&������8������8�U����Q��w�
�܃G�E�;��3SlṌ�+�"H���v�8�a:�~�Z���a5!/ܸKp�S�bv��9f�l�馗k��&���_��XT!�J�?emIY����M��3=�'	xj�7(>��֖�i�E��%$r7e;�������7�n�@��7=�]��9����L+�~�!x������� �iWW�:U,��p���V��_Zǣ!��u+\H�Œ�L6�<lT���7V֜�ap�����M �hp��B����#欲pA��uf�����0*�rFA�j��g�ccR��<C��K(�UP'�%G@q�)��n��W�3��;"�u�aW�3��5�m-EH	O�GqJ���<3/p8VT+�9�Ha=��!�U Ŗ,J��x�K���G���QAyj����[�yg)�"��y�M�(ͬ���8�;u�Q�Pt��o1a�X7��r�z�񔘦�ϣK�Lup'^m�~�S�N�S��N��M�ȓ#>�x�
�q�Q�ԕ���n��	Nt�fcB��1�	�p%�KD�W�.)�� 0G>S?\�nZQ�]���'J��GIǸ�ɰ.ó-���G@o���^O+�+�@onc�%��\��045a�=M���m�"� 0����^���0 ��\N��:w[��|��p���uw�qm��P�N�Tfc��v�XO�,G ��;�A��@R�d��l���>O��+��/�v#M��S �0VE�N�K�=������E"k	���i�-��\uQ�����݃u��Ǎ��~��G��G:��V;��t��ݻB$�%��JU-�.o����D`$6$z�����K'��{��T{d����,�Bq�4p@B�*�;��{�S&}V�R�%��zr\f��N��c/�B�T9�>�"|�PY���pD�BE�˾�ʔ��V'��`��z��Z1��V��`�B��V�u��Q;�3h���M~��V&3��d	��Y��[Ԝ�Vp�h� �a��9��-��O��*�9N��
��8 B�3���x��d����~A4��j�+-����kD�bx�|u��j�ZhkW�-Y٨������ǒ#�^����u����Yb�6k�/�w�Ls�ۓMo��h!h�p��כi �~kv�&�^4j��z~��y���rZˁ{�K�`Y��z��ن�&hl��(��%��+~��XO�
d	�=5e(����%��^QV=X풿�������7�������L�?X���V����e$8�'�e5�D�&���}��G�tWmW���q|@��s���:�@N�B�~5�f`���o'!uX�%t8f��������$��M��wk�n)z�
@U�C������ǧ$���k3#�B8�ۡ%Ċ[�eG�o��!�V�d��� ��9�ߡ1�R�0�!�~9�����1?�׋<��q��po%6�K�77�N��ȥ8���b��}wk�?Fm�l��v�Nv�
�{ބW�K�xŋ�8��`�*(�(�רo��79w4A��u���[V��ڳ/���ް2��r�Q=���T�'� Y�aI���,������aq���?ߒ�#��
/�-�5P�\/K;�<�����T�`pO�_v���L+�z����?�̬0ܕw�8Q���E�s�:G�	(��
n�Q۶��nT�i�c)2	�L�ȘbV�^|;���š�"%(R���[G���i�?�{Ǜ 4�b*�H%�R�˴:Y���/�.��+�	0�������:�\�փ�[��ڪ�G~aÍ����su�
�K{��I�!t��a`�W�P��}�]}|%>e�W�3*�=i�N��Gz@�Ʈɵ��|�d�[��4f�J�JR����)��ZzH!ΖnC��	}:�9-h�B��3��6W��A Yi�Lέ6=���4����_I�?8~9�Od@\o��ąD 5��@����˄��@f'�"=h�TXJ�X�r�5���o�؃Œ ʰP�V���N?�M���BsOs����M�-֡��uNi��tKb���#�klWo�@�E�6�#�vJzt:,�X-�;�-��Y�,��Y���G����P��zY�9t���8~��X�����i��2�Z � �����<�. ����{:킜�/�V>���
��159mw������N���Nr8h����F�K<�U6��F}�)�Y��O�
�����&!��������r0����ŭ!m��ȝEWQ軀*��#~�i��ƱyD����"������Ev�I�mUE[O�]��P�)	��BiBV�Opڻ=��M�� ���Tv$f�U��h���6H�!���Z�x�u�]5}��!n�Q��Jm}��U-�m���R����vk(!f8�{��y���D���[�ھ1�'`���K�	�V�ړl����O���Y���<�_&���	8W���&�Rǂξ{8=н�iā$�F�#���