��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V����hN=��a���)�硹<H��׮��`̼��D�g�;�mR�#rj��S��k@'�q�/�ha��pc�R�(��g�F�ו�����`d%D��G�qK�DW�+X���iv�O�O����9�t�0���`�<�F�2MGJ�g_Ю3����Na/��4-^}��ru1������>�9��& c�dN���(�lE#2���Ƣ��/�V!��"�2?�T���$��n��|�GR��
���y��������D|)|9���w����臧�S���J��wd&�Mi�5�HI���qm2y���GhՋh��g��� 4v��,���d�0��(�]���>&��O�ǭ+���t`��oƿ�F	E1�O�u��7`��%����i.��k�ϼ�U�l���}RoG��{��9�Kvd���0<@�m*���
�P����:A����n:��w
��G�K�Du'M	��~(2�'���;reE��OM��;�H�:���!"��b�񤈩�B���%�g��^k����2�{�E^���G&:0���^�o\�\��ٺ},uZ �b�m���T��8�@\� ���PsX��A�{d-ܽ�YYS�4�лz�")ʅk���l&��Cx��<0\�m7�5?�"sK(ȋ8٣��M��^/2�HbM�+����9?��H�oRi9�0}-�ҝ��Jv��k�p[�ZF<�L��\��p�W��[�[��+2��㭰�c��r?�a��+�ë��Mzƃ�y��S��r$�Ah�N].��=K���`J��s���Bsc��(@�/�Ct����~��Wm�}g�,�n2������C�ˆ�w��bV�W��aǾē����{`���i��.�'\��Q��>�J��>q�A�MO�R s��l�5a�7%b�\�? �ȕܪ�i�w4�j~�݁��t
��z�������!���է���Oz�+�d��z�}I�/	�/bE5���]�,�zO�׾p��\sy�P��j���@�=	AF2>�h�_GL�&�c
����-BJ������P���~��s���!> ��?a���T�q/߫J�qf�8�H���sr�+n�"y\���μ��+�b� ���qf8�oC�~&�@8i��ڂ=��Ǡ�Oz�e>�;k����i���6*�5�XS��̟��5g���cb���}u��Z }¼3y��|��"e-�f��Qš�m�$Ͻ�V�dz���uj��=c����j��t�R��B}II*�jk�#�O��Nm5��w�|P�x��cy�Đ�NX�,T&��!�e��Q���dR�,��L����dREQ$�0�����6�d���Vr��t%W�j�m�.cLV�xO��36���TE�y��3Y=���/)D��.�,��~q��TM�� S`o�NV`�����S����uY:TEh Zi���vq�1H*&��<:ιh	���g��Kư;v�'��s���Ψ�u���='���\Ρ��xߊA�GK�56�`8�`Ԯ��v�ǟ��3ޔ����E_�x��"�uU�(L�ǁ}�I{²<��:������(6ņӔ:��Kk��z�w^�zS�Ӥ99����gW��jS�`���is-��x����s/:?�*5��PZ�ޫ�\� ��l�^�F���aP35�Urz���`�Ē�K�����!�F��WVx�+�T`;�4�]�fI�$�˗Y��- �ݓ���'}:,Vd�`&���w���s}F5qJD��]���,��)&7m޶�aݼ) �m�ȥI����S��v�5������HY�UH��h8_xa��(�ߗt�J3[Ć�q.@I�n�M{����g�ca���|8&)�.g�	�����g�
!k��/�$���풀ԿGa������O�BI�[�jf�,@�qo���Q8��%�a]�N馇&7Q7X�o��@���c���1W��F��`�(�R	��\o�s��ޒIV�����6�&�7-/֕����d�^��K|��~`����e��M�8�V��1�/W|R��5}O�6:�8�n���ٯeqK/��3&7%�b��_��-�cg.��0�џI�aNW�
�'ξ����� �D^V1R�·pJ+c~ES2�#p�3�1�b��}P�������'yC!У��,E����f�-���]��G7Yw)M� x�r��V����I��<�u���\%װ[�Fs���xp���:C-*y����LC�/�X���W�����1���!)Gc�	m+�B�JX' ��"�d�ja��%�4���YgNKVy��)tR��J�><☺��0�8��6�&sN.ӡ~Wv"14pM+�^%#���ׄ���FaoK�β=��}����a�5��9k�a�_�Q���ڮ�S��Lze�+%>'č8�hv ΊW崣{�-�ċw����"9�J���2��s8�?�FZ2/�g�5�� wh�C�u�b�۶���:�uF]�%��kE�k^��F�~n���Χ0����H��Y��8��ة�M�߇N��͚�·��@Ty�7�+�����>�������0q�9M��Ma����4�����Ѓ����f����#����c�%���ǔ�"��3�^�>Q3į�pX n+�_e�l
�L|��_�Np`,q1�]/���;�g�b�(��i��H���'�9*.'ɾ7k5N%"[�\%�3yH	���0!��g�E�D�m@
�ۣgp��{��-��8�
<��w���m�ߛ����ړ��8[�o��}N���kU�Qw��tX;�|!�4EY�GīYn��2�O1�X�	�ΊA�R�NE�K�%>���>��6x��Ӻ*��
�IM
��9�c5)bHխC���]xkk�iyg�;?!V�|'�|U�oi�~���V���p ���4-ȍ[l/r�$6&�a@���>~_��L��7Po!��+!��w�[9˧�M{�MD�) #h��h�[��0�?������4��O�Ά3I��$����\�v�hÂ��#����I�P��>�5�z��Co��Rq׿��+�Avm�sǹ4!�u=L$�g��Gb�\�w5@"kg�-����(Ŀ�pM����y������*�)aK��T.r.:-^ܔ�D�𞨞���Z��V���|����!��-�1{�sKE ��U�uK[�)`�-pF�S�ҹ�|jeѕ�N�j�����/(?�Eѱi5T�~��}d�s\�P�tlQ7��of��b��42�ظ`���s� #4hZS����{y�?O��0�6��Y�J�2�S���OES�U�q�����W��7[SS���>�m��d����QU�Q�*�	(��ԓ|����<�? ��7MX>�m֖1�ި��`Q������N����®,�9^.�����f ^��W���#�/#��w��q8#/X�!�m��b��O֞Z�x���#v=�`$�.����H@@����^UR0fڏ�#�3Xg���a�|9�{��Go�. |E֏1�f�� P�>/ԇ�K`��d���F�C@�m#�ox,��{q����`��9Q�qzA��@���3��h{��1��/���X�b�@��>�n^�6�6#��0\����,�:��"�Ⲯ�
M"%
�I�NB�lq���,b�Ŏ�K��u�k��Y4s�ժ*E.����V��a)UHj:Hw�"��*o#/�8�NG�%�gkԋ���w�LŬ?2�ߥI���U F^�Rl�э�^Wq�fL؋��?��C���RaV�)
�-h|�SY��1A�
H�P�Ͽ�<�V�)^[b)��K��J���1��f:�~\Q��wӃkl(]�����ᐾ@�&��y��t�t�%l����G,���T�ۑjߪ�?ݐCϣ��L���z%������T<���j*�X%,
LK���@�
��3q{��d��ԏ%���1�s�4?���u�:��@+�3c�`N�L�4�<��3�a7kc0�ǩ����.soG����� ����3�G���&�"�ط
[�Q���|��=�v�Z��L��;D�/����$2���n�+��6j�E��&��� �bf��
uE��w�KT�[;�G��:I�U�����ǘJ'-�:�\}eVݙ��� #����b�>
�4fy�$9���HWw��Ԣap��~?���b�w��`�Tv�w�̬w����]���]I;��pR�� >��/*�D�$GY˅�5O�z�@�y� �*;��1��4�P�-�(�Y�@M�vW[}��4g���o�D����"�M��`Qk�A�S`��0 ��{�t�D�21���Y�\��6ἒs��"���=#�A�� V*)��ǱE�^�Ǻ#d��u�Q4�7?̦��
���G���[ o6dP�&�Gf#Hi�볭m�152�	A3m�/�C{�(wJ�;�諭�-�:�t��hwcuDЧ�߬VF7���<Ŀ`[<>d�y�8�i}{L��v���a����hz<g�Mt��T�eH�k�Mm���dR����@�����RӀ�Yo$�R��SB��LW��o`T?��W������ƾ��A3��S����	�p�L.�$�1b�!_��	�Ɗ�ș4(��1���́^ȸ&�fmY��"��5�z�նnE�`��k�}�����}P�+�g���P�)+S�F�W2�u�-�S��=Υ����M��� B"�SG,Y����_�.!V(Cdh��=� n�����'�s�X�H�-�Q��F���q����;,�o<.Ϳ�l1	ds�E�3���Xk�"�������F� >���p|C��������3/�)�U�&�7��|f}�y��=��+2nS`���@�u��JK����d8���I*Г谨��!x�Z>�썐�k�d�o�O�sC�LS����P��m9���nU�W]�l��4O��G4i�������=�Q�����ve�*G	��WNN\d+����t����G)��t�Αtϗ"��"�a����]j{U�0+?�9$�،CֶP�\��`��^���7��jB
�W���x��&0R�l^�15f�Q����{����� � ٳ�|}b����ۆ`g��M����!����[�Υ�K����>�F�@z���n{=���#�~P�1��oZ�)��_����m�����C[L}�}�(IrwJo˗3_Y��+��9���2KRx&(��U��p�o��-�Z���^���1 ��
�9����$��b��I�f4��3A犈)��֯��[U*2`� ��8"��4B\�Q�._F.�>�iu�HJ��=gD�,�#�4R�PLz�֎���I;��}zl2��i���̱H<J'��`���Z0#��P*8�|V�����]h �v?P�%��ⓖB}w|�
S�'���1���P�tL�-.��D��/���&�I	�����p�'�V6��Z:��(9�񳖥���iO{bܤ[�	�nZ��t\�J�1�:���}[̀�O�����F��K���D�7�4K�V�Z+{Jt��S>A5'�Ulw3\]G�Ɂ9�����x�V�=�(��y���O�Uru����g8��~BM�.�7�����7�]�L�(d��y�E�*��Õ��|�����~`)׏�����^��Bӝ"���eZvx=���I��_�F�{���2횎ǒ���077�0@��o�ʔ�y��q��y��\<!��F�)1��l��b��>I�#8U� f�x!X�[�4}IA������o\��K��cƦ6E5�1ohu,% �[~�5�N���#�?��fce���4��$ ۞l���w�J60m���Sn���	�އ +�X}�K�2�l��(&�&�lL^���j����M��4��`���/��C2b9]w����	C����������j�7�� �+���Fy)a�T%m�~�&�A_���8x!_b@
��?�����5�ZU���#�9�v��JP������dqO��[��Z�-�6ȋ��@�&��_e�,#��&F�:)�@.y�H\��XxO���!��3�'o�R�׈u �Uz�̢.�A�z��5�-�4�}�`��8� �u���A�ֲC(�[���mn�O��1<��f�������JnR�w�7����vI�����Z���OS-���[�7qH��=(�a��2�?z���75��B��*9-�<�@�0��wt>���
mSȯ��5�Ou�e޶CPρ�tI;/�ly_�R�6M��j�"�OE	l���h��~H��nuS�q3Vm���W�%��<H��A���'9)D���(M�urcT��4 o�6�3YZ&��K���9�����xa���{\���TrV7��S��e�JJ'�!���9��1*;Z�u��*�&���2���o�g������\һ��E؝�0J��7x����������Q2�'�E��d`0�M�������3z�4V�4����fZ{s�Nޕ��7U�R��76�W����
|��Ы�fH�S�QM��lY�] ���}yu�����~�I�k����.�(e�������K(@��%jC������F�6?p�*��g>��ci���O5N����rL�ϕ86�!�#;~.8�f<Co-��QAu"�[S��������GJ�UF'vy�}���|@9޸�� �;�u��r�� .u��>��8�Ѕ�ʥ=�d��'�c�T��9��;d,=A��E��^B�n�ϻ@,q����&S� ���P�Q'���zq����	����{5���)2I�a�%����ʮ�ׇ��y����0���}�y�b�O:c�G��\�&�*w4�_WC������O�n0��l�������;݅[��J��k�Y�sC��q���&F�A�ۧஈ���;4p�	��_����s�g�����%@o�Ig�A��YG0�k/vY��4���F�݊*(�Z[l�I�K�_�~��]w������c�M%�vJ��m[X��^o~j��$�([t@R~��z�v�j�k)%����&/<��i���jӴ�4���<ȼ��u]{�
�U���YpΊ��I�o�Il{���p�� ����ع|ǥ��n�O��;��t��- 
��Rs�@��&ɳ����<��@�l$2F�9�]h�[�*���(K*��T�Y�#{��K���I���u>��1Q@��6��v�Z����x�u(�#�n2r��<�E��Ҋ� 
�bЮ������)��~�[���c\#28@����ͩ�Z��+Hj���~�HJ�+��A%�SZ�Z�g�]m��ػ"ۗu� ܯ�H}�+�E'����O�[Vg3�rB󐻛L9��/E�`�y�rX=J<w4#;G��Oʭq�3���+��Mk����D;P����&�*��s���ܺ�������bL���C��̣K��}:��~�\�~��-2m�1R��QiC�K�b�W~�����{ 㥔�n��Y��<����h�d��+�|ʌ�p�?�g��_���G�x�`�Eԟ�-VV��ջ�G��A��mC� жt�rL!+	(�5�}w[�� �����ԭ�����繂�K��J;�K�����ZN��<75�w0Vm�W"�vպ"p���34O�Z7�b��C~sCȤ2�W�+�ۑ~H�B�p�&7��8c�$�ڤ#�m�X�D�F������b�{X�7K�oW�'É�E��i���@�π�~v"h
O�8Ҹ�����v7+��$�����jS�N���^��`g>	%O�n(!��4�cwX��	rs����7�J��:�arE�Zc��]U3��|�l)���ܫ5h(�FC����m��6�#< �V��E�j5�y��^�|�.@ԹR��9�ŋ���0����Ӝ,�S���tlڱ��!����4'��L�u�D�r�S�5�˝�~{�~ş҆�`�� ��p�����9��6_1"mӃH��r��>�l�rQ���١�Q֚�8B�܆E��7��;ºL���D�T���Ϛ�K�%N��&buO�0�{����{�qź��y�����E�J�A_V���F����#-��Ч�!BC�:�B3�����s�ix�������a��t���Z.$���˓����o�b~�5�6�;�*%b�r_�!�}d�	���zCÉ��NsX�ޏ�9�N�P�t+*�$�F�<X�"��2$��y诘4��E�yp�(�v�O�����=��H�aCK<����T����g�\ɡ��(C�B�r���-����h��`���s<1�/�h��G淈$@�/�T��g�"W�4O��`�v�g�7�l�X�OԼkKJ�����y���{:�,u�z</��s�6~����]g�j�6b�Ѣ�'��>cG��>D�ؖ)�!Y������k s��*���q�}�9��w�UX���=郲>A������y���E�:���%*����C�1���弉�Et�_$�]�&�mſW�n1�	*w�~��~� �d����)F�N_���f��jo�a�R\[���hbJ�M���FW[0Ƽ���010�,O�w�L�P�9���W	y*ĝ��L���+X��ʩ���U��96�	��u���g`Лo|�Jr�q�1����c�����H��@;f�L���pҝ�vWu���E"�z�bUʐn��P��r��c��Q��a_R���=�,�
��ܾ�"�Y">//k����yq��?�:���Q��E_����L���n*����</$2�v�
�	��T)�l�`U/�K�{p���򒙆��r�pCU!�b#���sE�y��0�_�@h+����?ð`Nc�!,a�!<�4[���-w��3��[�EN�l�Qh���d�#�ӏV�'$��ɠ��؀���ϝ�����?��~����Og�F�՝��=c0Y9��=zJE!r����.d�|�b��a��(�6n�a�����cM�Kg2�n.����ƛ�&F�0T]E���Y$�&k�%9����Qd�K�|�lVd"&�Z��_<��%��0� �M�Mʗ/�y��!�OH��J&���{��k��Y�.�T��"��9U:R�@I[)N����06�� 4x�]���7�r:�"Rt#��w6���C=<�傴�)��)q��G�%����؆�K�l��b>&�FK��O<�v{�J��r��M�aK��du�KJ�$?`�y�l@Q	��%��8k��E��E����Q^B����1]��@�n��shi ��F�>	,$��D��Ea]����9���q����[�1jl9��3�`*�>L�ٷ���~i�ʄ
=uv��)s��;��[#	!&3Fp\�_�1���w�Z���H9��T����;�A
V���i�g���1�x��re�R���3J��L�7�xԸ@�T1�P��c�{N�NOKVC4k�5|��epd���[����@��]��������w�ę2��5��g]Þff�Δ�UX.�A�6%��݃&9�ZgaD�eP�c�z��^&�Vj���j�;B:v�rs�+�!��!���<�H��'$*� T��4t�IK:`W�h8|�Z����X� �a�9�6{DvtX7�?�ר��O���[��h����<���B��+D�
�[
	���ׄ�5��y��7,6�A��� vt��q��@�t����L4�����a�0�Y�';���;�D3dU����5�^&���y@��{�x�%�Ea[�6�[�UqB�#L}�v,�L�~�k)j9=�����G�:Va�*|��mE'{S����.CD�tgS�� �E������u��< �����%���p�,XbwK[��U���%0A*�h�c����{�]2X�jZ���!�O�K]�!��F��6�����z��=͵5��j�ʉ��3�PxRN�)����T6��%a�LU�������[R~_�9�`+���0�c��3�k.�]����Uj3ȅ��x���t���l}���t�? FC��Yq���4p��`k���y˸K&��Q�@�u�����J~tm�Q�8�����u�QȮb�\�<jq����/��Y�������E*T���L�ks �U�L�?�Ö�(:�yĽ0�G%�6#Dw���b�ߥu����=;v��/��(������}�����8�BW�t�mn�pΗAj*r���04�U	p�d���oZz���J�8FP�̤�b�w����*�<0��o(������g>���m&�% m�wٛ>�.�7}£�}&Y�����`� 3�n������.x�W���x�	����̂���!��%@{��9����G�4[�Մ?k#_gYޫj���ϓ�����X�Lɳ�cD��s1� HW���+4$c�ۃ^� ������+a�s�)�;y��$!��`�C�(sjX�v5�r�'�>�pG��P#m��p�)�x��m�b(x�nu����P�N2����#(��\/�Wf�?�Q)16�d%"q���k.D3[tG��)���?u �m���`>�EJ&��M�)�
lvehHé";���p=��S���+A��O�8�]]�� �07�m
��y��f�:o���K1ݭ��	��� 8�!BR�C�� ������}�PE��`ɉ��qrg#��Fm5���X�{���a�R�T����V��2����Ճ�)Q>����y�i���B�,���Ǳ���WPc�B�4�;�_��k�+�	�|�4�E�{���J�Ѩd��C�ݭ��Y�
�@�\|1�g�kp�+ï�q� B?�y�L�ܷ��`���N�A��B�D���Q4��G'�v��_	f6�Z�+�Ľ�ȀCu�:���(��X�x.�}ϼE!&���̅�[�b�(����Aݢ���g`���G��qT��WPh�+���(��/�b�1M�&Va��~�z��S*4i�RQ� Jh��do��wfJ-���͉�S_������w|�<�"U4�oPz�#Y�uy,�b���2�O�=���]�J��I.�J
���b@l'�ۆqqs�n�*��y����0��Y����P[Z�p,�?ZLY�.�����Y�`�ܪ����!�
ܸU~�8����x��`!�׻yO����L���r����E�E��s���,��+GS�0��Nm�H|;Ih��z)��������s9#VB]8q�+���f[�q�r��ts�<���
�K����aN��'�}+ty���&_���g�Eֺ4�Ò��0X{�|Ά��-Tp�g�g��!ߢ�P��BjF���$?m.�����o⹖ܥ>�*��S�5eQ~q��R��(�d��t�Yah�H���}:��ȩ�Z�D��:8݅q�@r���܍��%݁�u)TozҖ ���>>�r�^ ���%��1�g��ż�M6��78�|J`�Z��|��muC�ҏ��H�2Ɠ��o*���˖�ž��Gɖ#��k�\���������ZC�3�J�4��~�0p��
.	�ْ�=e�ƚBF��*w�6�eCrMr:�k��"��ŭ�F�p�@�!�Ϛ�U�	��[\&׍]t-a7Kdοu��t���U��ۜ���˗�Iv�e�:P�f���UL��՛;�ъ����n5�c¤���ba%7M<��g�al?D��4��{��/i\��A.+��5�N#W��]~�`r�o�8�C<�.�
�K��H��E{��	C��ѧ�[�D�/�5.��v4So6Gc�^�J�5��������[#�{�҂(2�	RF��� �;�A[�ѵ2�*���[W��ܳj�ڨ��b�w�g�+~z"�-	�=&���;	*u?�Њ�j���8�M*�3f�-D�p�X�����.�EUK�B��xƓ �R\Q��|�g>��cUKj����$�zJ+��*K�Α��`�)fm��Ż�T�N�`�>�ȶ��}kQ�I�z�!�U��kq>Nk���\n�o�tsQ-��w��.E5�PP�YB�u���X�yY�7wy�^��_g��/���C�YŻ����	6�G�d;���C�K�W?��"zE��sX�> �&�#�� ������V�Oi��Jo��M��5;����8�s�\lƪ`�*��@��m^���&���q���.Ӡ@8���\��L8?RSX�wd����#]��IZ�
��5�])�����.9��'uS�����4�����=����H+rʷ�~p��R`�*�(o��Uʸ����NM;/{��~�;�p#�������Xۤ~w��"��hr٠ (F���0��OL-B��{�uF���R��ZJ/�U�Z�	������b��HjjX��'����tCe8����u��y ���vo2�Q#Ǚ��nf�2��u�_�Fu�����M�\1m��k�K'�9?�\n�2=怉{�
���EG�V�ʢ�����'���1���.c��#��x�� F���ߘq�ZC�>S�����Y�R���jzˢ3Εۥ ���F
.��P�>�NcetC3�d@ )3ǫiG�����������j��'�R��������ʷ����0Гi�wn$�AW&�� �~a��WI_a?�}��{�`\"؀۳L��5{Y߾�U'{��ɟ�$�L���_��G��=ls���|�;8��V�(C�#M�	wxj�jv�62��5��ҫ.�*���^ ����,HGP�Q_)z�X]������%y�2�6N}�h#k���?��(�M�c�[�f�ϸߤ�L2X�æ�O<��S	�4Ԁ���/;���⭓�\*���+�~�}�ܯ`]/ "�(��B3Lp��D�G~��{�W�0��R�q_�m����l�C��I78v�<��ܓ�!��$P����j~�?s�j���>:�<"���#�`/a�jB���̒M�䟇M.���$�6Ն�w.ժ��<՜V��D�6�|�x��<D�#̗�2�9	q�p����X�a=���ν�n,�Q+��ߧn�p0K& |�	�P;����l�����=�dd$@,,��L@E��+聨�;�ݼ�?>�.m���.Ю��i̯����v����O�lo�X���W^���ٺ�qF�V��Wkt@8;��g���8��ry<�a��$9�;Th"����=>�j���>Δ`L}���͕ӲVT��M*S�C�NfN�cse*������v���In0'?�v,\��-�CΔ*��6c��/�%�J��R�n�1^D�b��J�Tf�-�%���2WwY���K����ů���gԮ�����[£�,�7��q!4O�~j��[x��TA�O
��}c��F����@��Hqޝۢ~-s]o(��L�S�6��y���K/Z'���/\�Rw�٩���W���`-A�����C2�)?cL���S�d�r�v�ԝ��ҫ<�������:�s��;�9M�E�%o��ZM=���{�Ӝ�@�q�c�L8�hZ�LFHRVp͔D�%�Ǻk$�`���~W�n5�o�\���HAU�^�Ħ�L� <�'��^���i��/[�O�����UQ�zS=�L�c��+�pn��Eu�p��	�(h%��(�u"W���C�N$�+[�1�#��^)bLA��}(9�S��MzC��:����x��:v�(��o�� /��9�~C�lZ}�KRC>O/�ڙ���9|�r��|u�����r$������<�-�0ys�W�u����$q"V19���r�1���Q7�]<��K���� ��7C"�n�:���3�M��~u��Inq���X������܊uU�\Y�,�ڋ7�a��@(D�ä�5P���;A?sP�Z3G�/�����Kj�Ѣ�L������`��b�Z�c1"$�$���!a'���v$�H仼�H���U��P�������B�J^(#q��YF1�Q�r1�&����E��C
��}!�nZ��3Z#�\���E�58yݖ̘���������E�c��4԰H�P
�=�U(�Y6V�V��3���VR\eN"i�l��iN}J�I�G���	�-�v�x�'}�.%(=���10'��(a*���wӯ�Z��'dS3���_���E�:5d�(T89%�	z{l���S�O�B�I��,^;�#��)o��کa���$�Yo�$�L�M��ap��t=��Y�c�%�y4�|�Φ�XGcj�@�Z��j#����P(3��A8�R�#���{����kmN�Y?�	
����D3N�:&��A�[�&c����[804D�R���Ny�Q���������.����4/�{�6#����5�x}���Q]���2�O�£�Y���.�����5�jD��=%�80��S~M�}��Y0��8h(�Y��=ڿ~�@'!6=s��D�9j�q��~{�
�RjR�����y���v�����z6���_̓�ʕY��|:�k�`�*���S�W���:�fF�~�Yh~��yT�>�d*���.�`K�V���bGw��
ƇDy�/m2s���/b�g�(�����cy�MV�`r�4k�6/��6�$�H��)(`�Qt���M'	�̓��SE���Pv�훏Uo��'|/�aF�FU�gby�d0S����eW��PZ)�_�l+Ԉ�q�]���+S���xA�8����BT)��Ⱦ�D�
r���wd\+k6M���I�v'��~�wĮ����a�<T�Pե;T;�e��b���6��=��^d �!��j2	����ޓ3���_�����ghG
�]�*Z�?����7��;�i�Oq���%�R����8~�K����Q�Oy�<?��xBa�If'oQ�Y �~
`�vC�x���E�oa�ޔ�g�CHI�5ν��5?H�>��ɂ�+ҍk��C-�qL�f�w�Z�`4zf3���u�iuU�jq]C���)l�;gd�Ѣ����C��GqmT�v��SQ��q�of�@��ޤg4ď��n��C��d�V��s-6z��� �J�<�q��~�i�FѨT漨�%�a��\T[kdR9��:���:�Ҝ�[��̄gT�#L7F�?�|�i�v�]S�;�W�1Cλج1�;:O������-�=��A�/>+SY�����: ����$ly�5�Q�H��I�o�����Y�e�$��y椩�����2����p��/�WK��sf��7K]��u%N�rBu�=cW���S�m9��:���~�u�o~$��0��������)渂��ɵ��]�|��F~as@3�ͫJ�*n�|��8�8��G� J��i�K{ݼ�a!M?�����O���bZ�2���1���~)?�6�s|���-&�] �u&�bx�p$wQl�)c�}����wZ,�lҏ�q��U-`]<���T&��к�奏���#3�ۅJ�̼�%�++�ld��k�S�O�+܁�����Y�]�a1���^#d��g�5�h�)a����n)\��0w
��}�j 7��;�g�e+�7<�8�.Q�Yk]�~$Щ�,����r����(��ߪ�~�ׄ��*>�@Ь�<�����B���z7��=�k�=N��yW+������»�Na���_3P��8/B3�~�1_�l��X�ne@!q�lh�&���"�����ް>Iz�k%�7��ҋ��z�Պ�J���TS��r����!�Tς�(�rҴL41�d�]���/8��;^}���:e���'d&2����n������w(q4�\n%b~� �@��_�N�0#F���b��to� �$��>�8_'˂؃���R��岵�s޸�V~��L�HY�ìNy9%ׁj�ZcU�슣u\2ˆh��XL�L����%���hR#�w��&'������\��uMZeHR�`bv,�돸�o��Jm0�`Sb{�DMb�@�#!X�����I�,��[vMy��Z���j�q���i����;$�����G?�*v \L�_�0�L|�V�G�����}��|���ǳ������|N[���������{�H�AK���!H���4�����y܌��8�`�ҬcWbб ��v���&�(����i|�0f� �#�}M�8D�0���k M]z���W_V��uzcUE�)�L)q�o����d��\�:;t�����s����&k��L|ٵ�r��[ß�I�J�v�Wܢ��I�Q��-�1�<:r���d��A�xL�'��e�A���(;+L�	��{d�9$��O
	��j�5�i�!����0�= ���Uݐ:"55�6��*������w��ȯ��-�|��I+2�K_�O�ط7�1RX�)��T��+�@��a,��Im��2�B�y.6�B��	gV������Y����}A����1{�����`i�������"ek%�	�)�M�V��9�@������=�׼2Bve�!�z��n��
7�}����8$���D�[u9�"J�kȢY��"4���̟��^�>��-Rd�g9�>�d �~)[>x1��a��N�0���јo�/��~`���#8.Q3�����_�?������Z�SuXJSU92��u٫߀É�/Iք����I'��i+A0ޛ����莜��\��ge��_#�I)Ƴ��<����S�b�tP[Yp
�;�������� ��_9���Q�\�O\��~�
��Na%�Q� ��8��Õ�a�M���f���Y]�GD,��歠��-�:��桠���������MJ�r9�\*�7�[�L_�2	������z:� ��J�]��H�#����&vQ�Y�B�BL�[���D�@���R��m�
��i_#.	�Љh6���!{���W�,�j|�X��a/�B�r���k��Nm�	�e�	&��|�Au>|�!w#}�}�;�ҳ-��=h�C�*�;�����ت��[�N�i����^=��f�:��\(�����g,��`�!Z�����'S�p��T"(���dp�HD�q�d�u.'Z�xsL��?lwH��U�`�G��"):�;��E���F�IP��{c�u7 D����?myz����g ĵ�T~�b�D�����7e>�u�f�|�M��Pq��$�7H��u�Y��gk�V`�������1�\��24%L��IX�刾|2MR?�k���&��D�)��o�
�r'�HY�qGH��q��Sb��!D����̐���j�m�H-jr,�껷�\�."�jI�n<M��Z�
�ϰ�%s���MC�է]�(�����g��Ȍ����L��+L��0!L#��q��m���z�1cGWd��ax�j��H�"A{;����1K�È���N;R9��:�U�]ᕎ�6i�c"٧�ALU����	!~C�G]���Vb�пxu�S]r��̡��Tԥ);�+ k~��n{�p��ʰm����$x`�@KƵtf�A �:q:����֤>�_-
����R~R�gi(��K_���F����3�A'���B��|O�Ip��ܾ�of{���;�"����;�Ʒ��2��I�_�跄X�^hf,�MXF(��G����=��=D��.���<�-M4i�1*���j��2�x�8ܾ�}v����B�dj��%8�85R��ݞtfN蠈�ů�AP��dc�KBF?m?��@����X�H���xbGl�%i�^�S���6�����B�W�'�n���/b��s5"\�,���G�f��պ�bT�k
��㘌�qI�jx��\}zyᖝ	��є���֢�O���|v�7j­�0#n'��d�7x��Qh�a~ 2�`Rl{�ڬ���Z�!�m[I�[�B�/ |\�p�� ִ�p���ƣV���b������!���XC��������1P��W������ټ�H8y`��yk`�<�d`-{K傺�y=hӸ_���'���.XG�*u)~�3��A޺�䇶
���F l9o=�Lc�x!�d4���&!�_�+E�Q�9)�+X��ߦ��!�`� Ea,m��Fq�|��<<�Oq�$�MBK!��c���������A���q�rΕ;�x�Sc)�r"/��%��7�em������\��F�[*�n:��1����y83��hgb���x]��R�jHkv�7��|�4�d����{���B#J�N?�`f_��:(|u�� ���Q
��M����u�#�(��.�9	���̉	Ԁ�%�)��S��䶽���:�R����Q_h�*囷��&W:��xo�Kdz;a��Tb�XYK+����� ���w�Ơ�3=�:	�N�u�g�@�L��V�?]{��>�o�h���^gm��'�"�zJu�(��j�0����\�J��K�Drg�rfA�����}	0�T�fuT�"��q9,#�/������y��)��`E2���*׾�w�kxB�u&��5x �
�e���b�P�C�+e�G�_5 ����H�pnd�{N{ �zё8�Zzo&��e0txUˡ��1�O�$��L�O���5~�j>�H���*���1ͭ�ݧ���E�}TN�#���te��M�%&��>����ݱlT�E��4�/U�gۚ��f�UDo8�\W�'��(
�W�w����}�u�P{3|���!��ѳk/q��E"唔��:I���6�O����c��w�7�CQ�2��hĄ0�~ĳ��=�f��wiv/�wC�����.�['Dv䞿R	b�t.Y�٪�y{����`\*�vT$Ծ�!;�I��x����-����uJ'��%xY�� @�A3��M�\So)���3�N�RKn�U7D����$�Iֶ����;ss��4���K9q����wp����IB0�#J���T��m�|�
v�1�
��S&@���^�yru�5�H�KεNu�iQ�Å��*Mux�3+
������L�WŇd򫲰�&��6t`½.~/��z�t֬��*@ԺUZ �U���=�Ĳ���(��`��a5��à��	��B8Cs�@i��_����L�-\��*-
�N��OP�"��_��w��G��!�Az���3y��c�9�c�Ұ�5�����=w2YQp+gCC��I�`GJP*�"dhwv��c��Z���|�R�!�R]��7ᗗ�ԝ�j�=SܖP���mSb�J��	���jd8c��IG���f$��5������_*���%F��N׫g~e
Zޜ]�$�hdbm�m�P��;�gΦ;-_�Aw��{M7k�E|�s�J�	hM�����@/ݹ��J^�'9���)<n��9ׄ;xGI���'��q�_���GN@�+LD�5��6�H�	��mڄ��#�M�h��= ��"�5O0�y>ŭ��-�?���ԁbh��h��D=	�({��-`h��w��q�n����$7��x�n7nP0��|�=����7�I٦�'~�G�F�D����]�c,���W�&���B3ġ�� p�e��%F.pz�o�����|^�c5w��{�˧^��ï���x�g.B�?�g�a|2jĢ��墆'��6�ԙ&H�,]���v�ܵ=�I7���6K=G���&?.w��]'%q����p���u��~�~����g�$1܉��=�Ļ ?��f�ڇ|3.�����n�����!7 ��O��M�.�c�R �G�ɗ%/�V�������ʭ��O�L(�uͭ�=�%�g��'b�d�WL��PAl`�DUvD��!��[���"�P���x��ܚ��+��(C�.�:v�g2�}�Y
9��n��v��+�ҳ���TR�
�乄7�̞���f ~R��1��X�$Bk[.wcy���'/uHҜ�����)g�+�&1�H�F5V�ph�ͨE��KN���ʖ�*����I	���l_���z}������o>���U��&�D��vF�k{bv'g�<q溋�K�|�����~xR��k�6x� ���!X�?����@�mX������mAee���_�Hp�`��d"�N�/Q�S�ii�+@ze���-�	��h!�pw�9����/���`��ّW��S)�KC �s�mPN���f������E�����Oc����A��q���N�����]�H�'ZS���7]���q��:c�4�А��F�6��A+���t��z�
��� ��S3'2�7��0YDV￫G��ze���ΙƼ38����_rd��0夂�����U-^+�B1�5��}V#����y��k��}��z:N���n�P�N�;�m��[:J2؎�󻁫���@^�m��K��a7�,�~R�����*<6�n<�E�-��+-�3~�\�qh+z��}d�<C�_<�*'�c$ˢ����$(�?�yw�Ն���ER�0�@s�t�$�JL�Z�n|[��u��L;{����B��Bw�>���LW�����?�buq��o뮩��lg5���(�j�w��̹���q�&M��
(�
�����kv��D�c��������gwc�*ƐH3/�W�ˡ���3��P(��DP#��:Y�@&�
�C%��ب�~m��!1FU4���s|�Sm%3���$37�7cG�te6�$}����^����+.\�7��<���~W%p��犿�=#7^�T���YGH�f�����'�.��'y��]�E��?���@�EIg�T2�����p�掅��WPsQmpn�#Ĩ\���W�p�8���<Y!�ъ�����D`�n�R!�_���E��1E������Yʜ��3��F+��ЭΔ���Y�5*o��Kq(�z����͆�t&r&z�}:w���+m`�=n�>��fvLJ����2'Y\��K�a �c�N��&턥��Y���x8�jq
^������m�vN��Ag�jl��ևިv�s�������P|��l���'ŗ)=
�aגes�3x�C������x�� I�S���oiΪ��Nq�=��<ZueL9��&'�Kq�ysiy=Xik#��b�(���t�r�8Pr�}ؖ_��gJ�7�u�,q��PC�3݈!u�v����&"@{�lh`ʸqr�T�d���7fV�r9��R��/A���
TbF��}���/�m�K����]3������Y������c���KV��?{�]:��������P�)�J�c���X�ԛ�s����Ʈ�e�a����64�{�>��MK�f9�(H!MپI�jI��~]=�d�q*�	n|�1�j�O������/{\ t1Ob>��M�Yk0��	��N�_�.W��eFa��@7o���!=�w�@�g����4^�͹Z�1�C����:����\sC�?;�=�f������ƾ\*T���(���*ʰLH�|������ɞ��\%P+�9����>���P�1���u���0zV��6�{ћ�+���h
�}�і�u�-�ZQ��OO�Z+pv/Ԯv_/�E��u��	`*��2aN����m�m�,��9���ڏ�`n�I+�>����5B���:�7��qn4{���� E��A����Y��l�]�]0ժ��8��܋*�)ش���<w����Y�P�`����F����ǖ��,�\�(%p�� p#�������S>g�(Z$F;�* �aO��<T�ù����sI�I�76-*���f�=���c�U-�.R�<�	hʍ���@��rS�e��̺1����1��i���:E!�9�y�������~�7h�����M;͏EZ�����P�m4g:#[6ȳJ蕊�T���WY�����
�ܫ[�v��Yq1�o���p��N�
�9�|����JZǜn·)�]CJN�}�b��2���IJ߅,(9>��[��̽�5Mq��yZϔW�N#D��DA|�t��$/�e!^���'���b�Z���j��+�YB��mͬ���f�@��8+wL�<�q��g)��ꃕ�x4/1�J(����.���h}r7xMfY�U�/}1̉k���'~C�D�a� *ܸ���Ȓwc<׃ <ڜ�ܯ|i��زD-�������7cT�9�N����rYEe��3��A���f?�AsU�K5�P.�c�Ǽ�T~�f"�u&��h'��R?�+�U�`N��fg�,u[�S+���ڞ����g}�ޭ�s��4FHdT��?�TD��5K%������_����6Z��"՘��DL(�`!��TXy�:Z����d5���L�� ��~��)WQ�5�}�:ko}f�G��PFݪ�b�gQ���Q��&�V7u<w��0%d����i�/�Lj���ᘪ9p��^me���Mc�#���sh�����A_���:���}����F�Oni��'�^�j_��%5��8��Ii)DZ:����#���e�\I�BM?��ธ�B 8��3R���,eʹ:< a�Kl���K�!�8��Ϭ�!s�Y�H�3k}��'��H�]
B٥+�֎�뷊�O��T�ت�[��(w�s|� /8�s�c��g1�����@��X��K��yFq8�tcDՊn�ŗmÌ�nt�r���`"p�bH�!���`�z�Uϡ�O�J��Ζ�H]��6W���$2�㏚1
���32�u��p��S�)���ď�O?�����{A	��D�89�8�S��]_	<��Y�r�TpY�ް�����p��%?��#{���|X��t4pm]a���"Ph����S���-R���)�,شDi�
����?�<[���4�p`n� i�����홠�������}I�%aنA9I���Vk�^{@e����ѧ�+jW�e׊V���nM��r19�kG(����B)�<�Q0����Z����/���-}�m��8s�%_N�S~}�H�	�c�n���h�x�Ox(]d������
