��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V��wg��+��1�0��"װ��_�����/$j\�4�eWL}�:�Ԕ��P���	Ȉ�P.#�/;�b����j;li��(�(�^n� ��q&�w����+�a���\��J ?#�r�xtܩ��3�}F(P��G�2�H�r5�$�2FQK��@���I\�������ސ͇�,�-�'"U��b�'�(	�s����C-dO#[H��.�N��|�9�>���sĐn��K�A��?N�������Y�j��3�0�!��߽�p�a�7��D�a��Q*c�B�(Ӣ�K҈�7��wB[�U������Gz���\\I�Fܩl�0R�T��-c�
�A+�K��j��FD�E�82ǣ��}�a��IM����lZH�am���׹�D룺�Q�9�6�g�(�p/}J���y�eV�u���\1<˛ʤB�+[v\a��t�_�Wե��g^cu�����R0D�R۽���6�D0R#4`�����_���8�٤(ߟe@�b��K��o~�t*�0H���7�ġ��9-D�e����3#�'��?�����'9a�'<����R8t6�U�}�:{�s�� ��p�[�n@�(^���s��|hr�&�kv�Jv�h#
+u� �d�>\�
U#�H�c�3c/�����^c��kO���􋁹�O=��6fw9���X�ˀ���3F����尗Ư�]\�$7�K��$WR����'�8D`t-�C�*)C� <��x̫,��_�
�9��Шq��qA�
R�eOB#�U�e?�Oҹ)�U�i)��#�Ʊ���K�6�Mr�4�>����5�#D��?��Z	P5�W�8��u��L��#��.&�u�(L@K�L����zο>f8�cq���W������n�{�X��;�Kv=�"��di;�n+�Ѕ�5d�F�I���,�iB-�|��[�\��C��1�R�ܴ�Y1%��RNdN�`�4`}^X1�k�W��H�e��!����G�r��IQ��8(DoK\�f�A���~��1��6��7�X��P�H�U����CX)��U��gk1�@}����IŅ�k%ׄ��8�M���E󔎫��L�A���1P[nbqt���k��cO�q�4G�ى�dW��y�����T���"\�h�Q�h����p���:�>�=��ql�ȕ��~����`�(l9̩-�����}�xpi��jA��t�w0}y�2��3�2�~%&�X�1Jy��y'�FC�+���3��*Ca� �X(��yc�D5�j@j�J�v�ы|�\�bM���^n�b4j�1��J�,��c`��\�w�D�B���p`4�R%ӣ�C�X|jqS��pE>��:UG(�~�~A'!0$Ղ�M�{���	��q��RWC�ʓc���Pl�9�C�����PE��z��k3�j�j����K�]��nN��_�t_�n�}�w�-�M�ڶ�%�Z��	&�G���Bwz��	i����P)���~(�zPZ����3�(-�2����PK/��+[�j�໵^
����v�xcY�x�2d}g�9�pYr5m����h�2�V�Sxu����6�X��iGm>[WF��V^DLF$�j�ޤ��o]!4�qm���-eז6�K�;S�*�xf���F.�8=ABK��Ea�!p!�y�c�"�#&�N�);8��
���K��l�`��^�ެϽ����C�N�z�����O��H�P��Ks����A�)p�z��R��� +��2�;��ۧE��J����1C�-���b�]�5&�T�8�F�Z(S�!V�:��%�.�^�O��������h���-�#Y8BϿ���ʿ
��&�)e�m�����o+;*i���ڨ�G���$��ڷ1(�n5�V�
*��Yc�]��L׊Dt_\��>~��w��k��Jv��!�����P�LH���	�%td�2��|z�F�*f^N��J&��W7��,7M�3������Z)�У��O8}���/
�
�,�k۽��K�A�(K~�8�m��q:u��W Z�`���A�=�2�n6}�R�Sia����~���6�D���,�QD`u���H�$EV�&\e�2	u9Z��+�[��G�%�kkǗ�����(N��!�L'��<i���t�!�hX�=�m�Z/�Wl�`�,�`��ԩs2��k'���y�����@ Q���IO���]YS�M��=����^�d�
�?�h1f��G��hJՠ��$r�j�/.���%�[|'lr���eKn}��3y�n9� ���&���];2B/�S�8E�1IN$�x����H0���w+^ߧn(��u�����|�<��w�v(#�(�
�G�3��,�t��ڜ��SO�~U;�2Z$���6@�p�`�9AY���Ŷ~e=:"&3��l�f7�'N��.�Q{� �:7%�8��eO=0���R7�}1���"]�V�5,Y���4C�F�6_��I;�g�:	w��1��06�|fn�	��I�+5*� X�k]6U�N�s-�K=��&����]���>�J����3(H�]���������0�ϟi@g1+	�}qz�T���.2z��u���DF	{��&���{���,a�"8��PSLe\���A���g_�5]��3h�F�7�粌3I�v�{�Ftr�ܭL��Y�z��c��_����}�����L$+���(�9�p|hG�R2L�/)4�qB�s$t�n�7R�B��r QsU�;�����<vouaSq�8lXOs[O��,�W��A��EF'7�96�a��HG��_7j4�%Kի8p\�*�A�F�#�H>��B�2��a"4W�2��r��Z�S�6�H�d0lf�?�\YJ~閜�Ց4U�@���O��#W�'�3oU$��x�'*#Q�C����FmJ����Z���i��a�HQ\4wnb������w}��oi�i�`}#(�߫�ZҾ��2�� �������ϱ$j�
%��o�JZ�8�V/���ns�9����O����}b��ʅ 8�]��_9<�aD�'uX��
;�G�����P��7��xC�$ �K��� �m���X�`�3[ɓJ~�*_Ĺ �v���{W��b��7E�7Ne`� �`�;�N���z��Ny�z�$�A���V���N�X�?�H @u��6-����z��I�ӡ���v6�w��������E� Ȉ���x*�h�3f �#g
��ϝ�W釸/��u��U��s9������'�ȴt��*��iùdIkl#���DY� ��\6W��䶵
ɛ���\c�a�����@���F�O&4����s �)�vx|�x$\��Fk�
���y-����W�O�8�)x�ݽ� �s���Y��xl'd��"
�hW���H&���`���C3�E���GtΩ�w.�B����@M�"?�eڵC�/ �"����OF
|�pX^��p}��LU�����;M j���H�O��� �KQ�긨Lw����*H/�Z��"
��ʇI?�#[��mȘ��.�������ut�=���sɸ�[�7H:���:��)L&O��!�����` ����9rV#��s��Pk�A<��	$m��$��.������۸�������.d\�dos�Ej*��jni�o�R�6{�?6����z��kx���;�$��
�l�fB'�,�Bu�DT��)C�-^��Y���e����c.�ӆ�]���-3�/gG��Y{/y�QG��%�[�Xcٙ��.����)�qT��?�;�Z��+
p�G/�v3�dD]��_��+��Xw5��Uvb�7Z�Ek5.w>2��p�e{�o@c�Y��A`�F��b	�o����nG��E�t���� f�
�w���Cg��U�KX6ƌ0����&�7iHX��?*������F�Q�N��b\-�3I��P���^U�8�"����<����&A:�����ү�oy��	A���/J>%��u�iP�D��#]% .�R� �ska����{rY�V��d����r���^=��k��AN�s�����-͏��{�e��L�S��!U�t�R��������-��x���O�',+��y�ү��H"��^L�Dcl�MP����u�)�+����D#��tZp�</޳���뙈�O�\݋�D����i�#���\�D}��Đ�ȣ�����K�I�M��>F-;�9k7m$e���ݒA�F���e��q%���vo�Rr���
|{��
rja|�EXxE��y�+(��h�e��Qn����Y�!]M=C��a�޼��жQֳ&.�z�6��o=�=�n���c�<l9����L!��%f�̷yt���f]�Y6�[�/Y��z�y�Rϳ|km�[�D[�6��kv�DG2�OG�;V%�4 w��v�`R�����p���
��?��	��T���}!$wm�V�Q{�i.�ځCZ����ݒFb��m ٣��/ƂL�����]0�)Ԝ���y��M��GV��Vt���n� u�{wjT9���vQ6��`��b �2Ա[���WsY�#��jc�d�b�2	G
�,o�ckaZI#KK�%�/t� ��΀M$~9�=�c���-���-5H��5��jʂ�J8�
6ɯ�$�_�������q�^�N�d_���)�%��������^�W0���&��"֜?�&��9�+�1>@Ɔ貑)�������