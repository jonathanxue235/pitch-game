��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V����hN=��a���)�硹<H��׮��`̼��D�g�;�mR�#rj��S��k@'�q�/�ha��pc�R�(��g�F�ו�����`d%D��G�qK�DW�+X���iv�O�O����9�t�0���`�<�F�2MGJ�g_Ю3����Na/��4-^}��ru1������>�9��& c�dN���(�lE#���{��5[{��X��������dD�O��������B|6�V�?S�M:�������!�tU'��]8 ��<Ŧg���f�-^�,�_��l};�-��['Ͷu��Ă��A��u?�Ƚ��.���|c��W~kG��G���Y��N�����n��α0�#�yY>F?%z�W=��q���Z�������M�N��83t�RF�%����b��]��<pG��+����X��I'z2�:R�5���6�'��K�3�)��9�#��PO\G�ڲTs�����E��7��[�h�]�XĤ�x3�-��&]-��j���8��	��CsY�cN��9:�J�V�_��`���M���� �"�N�!U���P�?��kV��������	�X�$�b�`������G�f���咅������.]�?G$N�����KJ�9OO��8(%b���

^��. ��c� �v6N���X�f�����)˸B"^���z�5�ً�;��jR{F�|Lַ�v�U�r�ų�c�x	���EhoP�A;���A��M�"i��.�-6��&�T��yj�G3m�!�����G��=�ölH��!w 7�8�ޙVa���g��%��)5ua��'�=�s�4�����5��Fe؇���B}e�ݢ���ʌ��'oU�
S�"�P&K+���ԅ/k���?���ĳ��#�)��Տ�����adj�v�����lЦ�L���;(�!�9�� ���N8E�{_,��U����!Bާ���[|ݺo�Q"�p}�X�Np���e �zS�+P���E=FV�������R � x��ĭ�T��|��m��;��4�8B)`�Pl�jL)�����>�w�0���8.)��9��2BT��(�=X�\Nt|Ӳ"Wn eG���)��������_�Dw��|'i���P�D�ΐ���Tr�Y٪�D��RI�y�B-!I�s"�襑\<h��u��wH-~��`��5� m�s�ɿZ�{D�"��cge�8}�,x%fo�¼��N@jQ?컓����kW��������C��da�,���ʰ8��3���,$+,�0kN�(?�b��@?�P��eB}�}dXi�X}�������vq�< �<+	�׆�*$�W��H=�r��H:LD<g^8��+H����2�%��im�?�,��)B0GsGS{}���u�ht�x�2.!��ӷS��8�h�DmFȽP��,(Ԭ����3iݪ�&&p�Dw	��b�Q,�O��[������~���z�Q�O
�>=���������@�'_4�q��7腝�s!�����i��?:m��M�C=8��&�EU���@G,���a�F(g�ڷP�T�)}U{>�n}_���Ã�?���⣉f�2Soa�� vd���5����D��kf��ږ�g2*������Q<�"�l���tpY�4U�����C��	�����qQ��ɶO`:��$������q���4�&����e�5�u�`�L��"�?�ϕj�!kz�T����ǲ��D�(rJ����7j��Q����{�����ʐ�VV�:ov�9J�A�>��6���q�<"F�W(�<��:Y[|ˎ�8�h820F��� ��|Mx�Vn�Ue�T1�veO��j�.:�F�U0�k*�wQ D�$l�t�ʣq]��+����91Ah�ڴ$ؼ��}`;0!���U5E�+2�Z�H��M�ʂreX��M����m��O��RiA	�y&��3��P~b���
 �a��?�1�1�W�_��?��㢉<�"U�*ᧄa�o=TSfI����Ōh�yҺ�K�����W+Ov��y���~��)��#%�FہA�=��iS<�	�I��P����S�T'�]>���=��i$��|�d
�Ѕ���d����1F��OW%�1S4�9��_���!?���m�PՑ���!���&#��&�зvt�`��
�*`�#�Dd�忖�rv�d��Xɩ��)�<�ѡ��Ⱦoz���#�@Q��^C	�f���]�]W�P~!�!
n�H���;�򕨄7��i�?��_���c��	mo,���c�&�7��A��|�YD4Q�}�ŭf5Ǐ2q��� �����Q���u��'��d񕫓8� V@t��J߫(m�s�Aa<��y��z�@�up�3ݝ=|eu8l�\�!qxsL�
�Z�S�LA�����V����p��`!*����$�L�[�Ջ��[�:��J8��kVx/� 'M}�H�0%��;�15��
�.�%������?��G���Nc���P�?c>o�S�1M�GC-��YJ�?�n�������zP���"?HXG�n h�
w����S�\���MG������?&�*=0V�@�8��#w�����zn��Y��~���f�`]�e����ǸY��+O�D�B�IJ��07
���`]u�v|.�u���ED�+|���/i����[�W��i�)j�No9Мv��9������F��
ۍ��&R����oV�+��k�nJ�衞����Ё2@a^��Z���$��VCNi��6�m�ت��z]�mަ���H��
�����KUT慄���,gl�}��Ԯ%�M�	ݖƓ�D^���mZl����<����!�{\�Sa��7��B��<���u�#sc�xB�[W<X���񞕆���B�;En� ���
{xMyeou�_�z���(�#m�e���0_ TF)Z�HL�_�4�U�!���Z
��������2mY�m-a�}�_����«$���YT���e�tX�GtFҢ��d����=a��ʛc�$��p(PuoJMha���wq�����kyȇ}ȳ��rb����7�X��J�F��׺���C��m(}oW��B�p����N��/�)�u�͢�>ә�[���=E��q]�b�y.,Tzح pE,��=�Jv�r�ê�7�z"N�.�����*n��:�JU$���BrYG�y��5���j����G��7�ve�4|�ϥ�`1�_�PWZ�ۨkVa� {ûe\:���.B�(��d�	'�d��C8q*�o[�Db���j�f�}�Ն�>#F迵o�v=3��e��iPA�����*|Ɂ_�B�	Zh�8��v�G6���Ȣ��N�l�m����m��I�]�$����O��:� [g������Z�WG�K2���)�X�q�q�C9��#�3��l���C'+�R"* �h j�C�ms����<��L��ܕ'$�PմN/C��[+��������g�yN�G�K�MWN^��%y"lj0Q���"��8Ti��Ʊ�C�j�pF^,�@?(�(��^���]�W�]�@���&�8���w���2uO�?ߪ�JX��1����,�.�]�ZF[6�E#;��7U"M'ʳ!K��8���ʮl�
<L���.� �3E�b�[Z�<Wh�R!SG��"���X�ࠝzgM�������SV(P�<J��g�T��s8�&d��w�H��4< �l~ww��q��,�0R�Y'�>�4I��RF j����h7�P�I85h���VϪMX�gB��>xb-�a�ɲ;����@)�8m��u�vܕ}���(�����%d�$㬃DV#�]h2�l�me��m[mZЉ��X'6��wR�H����?52�gy�`�B9��1��/�,�fVz��FN3�b.I���3������dL�W�0�hN���bKџ����+����[չ�����'����c w��}_�2ލ٩��To _��		�����` ��SQq�����+x��ci�����d�s K��RLͿAY��3��A`5�"E�_4B޻����J�y\�n�&��5l|���P�P�lǂ�Rq�?��6uM� �o�%J�n�+��ӏ|�)()V�at�f���zI}t�)�(H��tU!�u#��C�OV�( u7���@ywQI����R*�1��� o�m�b$,|�./���G}���}��y�^�$M��!I"w�Ĩ^8��!N��n3C� t�*,�ɚ�/v��{�]/İ�9�vH۱�$�)>#a�櫛�����!E�Y�['ΞU�M�0�=��Յ(�,LQt�׽�^v����y�@����K����~|��'
J�0Q��'׷M�Ú�`�chAt�*sV�(cBC�����ڼ3��e����_��/�O�-�07C|�1#)Ioz-\6�5B=�8�A�G��o`U�W�'����h$�_]E�a#!����`UL���i4�袤����c�V]����8a/���|y�_��-���@��E�J\��Wdע9���Q�b7���Z��Zwp�ߦ��T�i�^��>>�8�`pJ�gXQ�s�7��(C��}�ԏ��W�t��45WMje��bXwƕ$J�F����4`qK�mw��f�u���uIj�))N��m��IJ2}�)nA�jhJ�PE�l�����\��ZBM���mi0&#"dv��(X)5Ħ[0ҳa�P���S.��e^^q�O��2e��2|�\�$�f���fL6D�F�F��&�X&-�Ym/�<���-��i���C����&t)x�ޙz�4���(��P�~'߀5��u\�]ȧ @�%H���<bjT�f��d����5u���%��&���J5��n[��ߤ�3���i������\�j�_m�ّvl�3y�(�iH�k� ��q��O�.`^j����xw��Ueei֓ϴ.1��U@}$F(�v�F6������O�/������|�C��q�n��b��v��e� ��6ƽ�d3��}x5��6W�U�1r�d�.2.}�2o���w��êٟ܊M��Y���R~�3
���e�����,T4�	�7Z!���}��2���6�n��9*�<f�O�܃˅��/w��i7.zP�_�q��̀���[���5�����Ι:����\V���GY$�K��]���w���3;��������2�:��js���-�����;�F��VC#� ��ףV�)�]ܼr@��0a�{�@��y>>0����;lO���=g=6
�f�.`4ǺDq�ͽp�TX���9��h����n���'����&iQ���|�-���-���4o(T�b��4ኁ���k�-='�I�A�Fd��[e��z"�+/~3׬jn=�E��0���ʹż����9�4�o��ntζT,�!T}����D�6/�9�  ;�Q�2����>��V^oGܗ��ʝ��5�*2!�������7#9ܲ��碨Ã��	[����AJNe��k�&7�R�O@?d?�R*e��7�$�6�����؊����_ ���0�)\Yu�x�伕Ny0Y �+���Q�bxo���%)�$R(�fh�Mc7�$J\O<ppq��t���-�S���z�d}��j&j^�6?���f�=���$c�x�[J��-��n|��n(!^�1߁��iv��R��ǚSX$�y:�sy��HJ^�{��I)je8\d��%�����b���e�k�1V����$q�H�S�|U�`�Z46m.�i%hު�1�]|��b��_Q�O-�?�v-�����=��	��g�^����9 ��"Ym�Hdu
�Q$�+1hY�:	�Oہ���pǩ���ף�Գ��iD�K�=�姷)�Ί)��`�����ˣg�*�J��P��vk��
�y����w�c����ȫ����F$vka�.�*o�	��& +��Bg��ȵ3F��ze!������q93��w����]Uq��l��/��XKWw��5,�2�Y�.=�9�1G}�O�lkz��}]8XoT.�P��.J,F-WVk�cI�ٴ�8���p��n�Yl�,d~��,-l`%σ���*�J֟���h���ک�=���X��"����z����SK:�C ��7�4
��&-g��>�v�Q�c�繈N��e���(���oPһ�v�O��w�;��ܿU�JBT�2�¦kr�t��y��?���	�1��܉4q#9?_�@�1p� �Qn�@U��D��H�W'H(_~F�����hk�2luE ?	���h�ʥ"�=�eS�~|�pU-EZY�<~Ɵp�� �'�&��>�Ȗ��c���}��l0��fj8[I,u��bXSҙ���G�5���$V��㠯*�}��,�dϡR�� �O��'��ոA�[Sty/�dP������Jn��f ����r�15�\��\(��+�@j��)�ಥ.����]
���Y��#�t/�}��ot��^�������B����Z�h�X����9L�&��ЕsxpIB���E
�F6�/�٬�g����K�+y�p��x�M�A�X���	����,��޶-F��2�,:�8��Z�~Y�ǲ�{'�yZ5  Ǆ���N#L���1#�usO�tu ���Oھ�.x5���̚3%+[^�M��t�,�p�x�÷O6翳�PnwQ34��[��w��3R�
��
��X��
�\�e��D���hmU\�oL>��쉕KN*i�H=�h}�y[��\y��k����6A��[]�{C;uA�FԲN��W_�S�G?ش�O��G �U�R�RC��y���|����E)�UG0}���'�R`̡�KP ��k���8Ȣ=�#`��$�z��I���SP��w�b�L�]B"^tz�������妟ްфj�>�n�=,Fʗ8�r( p}���1 �q��-��>�Рw8���o<AKU���\CE�&��ř��|��I|Ý����_�7j9�����H�Z�"W�O�v,���bi�! m��ǎv�5���n�.��p�������;�	�1�㴟s�"�a%�a���Y�՞��.�w� ��B��G �XE��&�0\}9����W��\�PN���ME: �iT?��-ωwJ��C1�\�����7 4���"Nc�刁R	���iF�X$���w�8k^#�Nj$��g^�����Ema����Ru��M����������[J��rsR���F�8u>+O��Tl�*�#�iҠtFC1�UI��,��u9�-���c��>߁����V���e-���G��͊%n	X�ZM~S�+!�_�����[sj�PҔ	%n�?�Ed�P�߫?�q̑���� XT��:��ӂ�3��u4������E7����I|���zxS�+��8nH�����T��; �C����m�+5 {v`VD{�:Ak�&�#�!53���p���%���{>��NՖ}�V��/�-Tn6K�@�MB���Pa`'�׫�bcK^)�R&0h���ț��&i�ju�U��Ƃ�)�3��@6I��>�^�\��Ǫ����y�:<�wk�����e�i�!sC�P���>���])�,��NIaA�u�$qD��Ӧ�U��c�J�	uv~_�c��)<yu�'< ��4��s�%���ҳ��=��YH�i��?2��o~����N�0�t�����|��ٷ��3`�\sΦ9 �6�W�o\H#�)$:�mxՉ�v�Q���"u���S]�w=��z�6 �`)})�TX��wk�"�*B��=��L�Q'D���?���[:u�֛�-3p�&5�8W�#C�~ȅ\��~��q/���Ͱ�z�L��l�ÿ/-��.BRSq%����B�l8ca!su��d�=��]-?��HL��ɩ���C�e��R}��TdB����۳:!#"�6��\'̦�M�f��i�<��X���5����&��gE����6* ���~���$�w1Bj_ŚCX�v3���z�`�[?���]��f��������[Iex��BL���kϨwG�Ԭٕ��ĉ9�|�v�4�
��qa��~�Uԫ��rzy�GQ�7���>�f���*���1�ui�J:�-��}MLU6�~���C7I�`�*_ExX�?�T�c���\��NDh|�.�zAM���'l�f�A��I���Otz�AS�I�1�,	_�����tD3�#�{��Ns��f�r����4� ��;NG�]ݬ����b�ԙ�PB��!Z��`���F�VzO�?�;-���Vp�~jOT��4���6�o��[���.\8���'�G̲�xw��t"Zm�Vh,�u�u�b"���km�J�yO�A��LRˢEC��<��D�:��)��OAV���g/�Q.�'��XŎ4�M�b�ZR>���?�x�o�{�L�z��6��2�3��A�j9G�GL����߱=