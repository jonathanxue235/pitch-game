��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C��(b�g L�N�W/u�b|���@Aw�_��5����w��&�T�`x��i�>+�_^�u����V��0�d]����w�������x5?�\.�r�A�O�R�s�s�l������_���eδ���9��<k��lիK}����1��0�f�?j�	�l�֜�e�	1���U��s�:�$ɻbB��E�Slo�"�R��U-8�"�s�0�gr�=�*����Z~������ѣʫd !�k&�M�v�}��"�/�Hbʩyp�N��L�z����K��� ���4�p�:�X�ļ�0*�Р�"A%8������4@�+��}��Z���e�������Ƶ�r7�	�0aMj|1��2}[���\�E����E�x6S9��k�G�`CP��S�׊�E 0����g����q-�6����O稷�c�>�D���-��
($�5�
�K�DDy�v�]$K��ϊ�B��1 LhӸ}0������K0��_x�:�Ih/t��e��%t+ɽ�Ȏf6�bhu��;,<#�H:([8qr��,�����1Ȋ�H�Qp�s�f���y�`�a��:7���F���"7@���;��?��$(:1�O�[,J��\;��5)b�H�XzvK-/j|}g�?A�
|��J���@�?p����<�@����!kj<�M��f���<���G�\e_��4 �I��q��z�fw0���!С02�Ɯ�WH�<Ͷ���h�%�l�xU~#�-iM1�m��i�uy��Y5�*">?����	�*f���A���R�W;%g(���0����̮RG�@t+/���:��~�KRd*��SS��)��k.{�\S�9�|�24kW��8���!G�k�Īʊ��������5�WEa�8[��XfAJV���-LY�P�Z���W�0��rV+,��^��BI��w�6<X=����˹�4���U1Lr�b���%2��O���f��,�z�O�2�m�R���F	��Uْ0��`m���F�H(��W�*Є��K��%rĩ����z����^�wf2��J^	M�hZ����f�/�q2-��q�"�س�k�{L/qڡ��}	��}�4�y
��Ƥ��5,O)�����f�Â`�{�[b�ps�-H]
�R��Um~	̩��Ah��#R�EM���Q��/��Y/6����v-�8�^����v�q��m>��W��H���s7l�x�)`ĩOB�O�J6*$|��E����������Ts�x溔pN�7�#�XSP?] �����8�B�LȐ�{ӷP@ʘ�:K5e6��7۵�)���oN%���eg�ආ焯`ql6t�PKTf���wgI�2Nz2�n�Q��5���$�l�k�{f%E0�k�߃Z�h�
��7� �e��.�K��� =���42BO�7Y�c�H���e�e������['���#�U�џPd�m"@.E��k ���ٗ��r{B�-f 4^x��[��6�<����Z��펃O��%�����
?�~�sΩ_2_p^v� M"��,O9�}X1ZL�:���P�������:-Fĸ���s͸�߈�~��eҭa��]y�@��f��D0�L�l�kC��k�#�ɓ��oAFVyL��@&����0]_�� o�B7R�G&S��o �mv�A	�أo�Hć<b���70�_������%��de�ú��DL�6x���߯��]-?c[�ȑ-qF���ob������4hE>�:'��yo�e*�2��r:	{�x�E���(��fBg�T�X��1d>Fܗ���n�_���~>c�8�}	:���.�����\Gg9{�
U��W��`ᮬ�t�6pB���n �a�^J��K�U����A�ⳎC�6���;4�,��jG]swڈԋR��$R��uX ��x�_��񸉌ih��\��h��}�7�����ӆf�$IA�@w��6�+bk�WϾ}���w66E�S�_b.�_�Bĭ0V�1 +��|�j�%P�e�k=bG�F��&��ۓ�:����J���O/���~$X��f�㸏X>q<ɟa���p��	�$ix����~g;�����\%���j0 #����w�[.$�
C�6�[0�SO�A�K�'����#\�X�AY��D��oa�M׋���h݋�&��o���𼝳d���w(Zq&��E<Mu�=D^<�9.�ɲ;t��N����<�=���v��Ǡ۵��u��Prʹ��J�\̧ 4�
v���� &)P��7����_���/��9�3#��%�n3ot@����'������$�N!tobi0��Z�L3��K~�yg�}��s*�o�I۶��b�Ä6h���X��{O�
$��/�4��Ȥ����R|M���Ž�++���Zhg�Z�2�f~t��
��^�3>�Q��WR�oLdz]՛�������
6��1�f"_ef)����
~���a.�2���B'��8��
�3~5�8����Gr�Z�P��(�p0��CF�s�������:�ZlN-����b���.Np�{i�I�� ������F��`NT9�_@���
Wglc�r��Y;n�0����a�h^)�V��1�ר��k����g��!���[̒��_��=^�����]z��՜v�F)am�_�W
�)��B;�Y����fĩb�(��(ma��0&/t��^�Qrs�I���2�V��0N03��h��S�3�V���&KDu�u�f��������z�� "����\&��V��s��E���a
"r�� HP�m����Vk���ٯ幕S�B����GΧ�|[�+��O5�R�����-z�S��2��ι�b��J�F� ��
�_v�1�;�P��$�J��.>���Ŷ$���$�& o#\�by�Q��f�}�o�*�<B2w:���s�Zw�h����P!X�c�D�o����$�&I�=����w��g��=�W��uS�`,��>�Q�C�C5S�6�g1l�~���s��o����Q!(�)¨b$gw���?�0Y(K}\���iH5~'!��uH7�D��x�gVaH�>�2�nA:^W��9�l�\1���{��Sz_�B�x��H  r�$�1����!��u��g,�"+����,q��&M4w��@H�R�@��`{OL�;�t�ן���a��Gj����E��������i�O.��<S�w�1����De1DD4��,���q;qQ%Wӧ� �56�N���&�����e!��Ɍ��䎖I��-)�(�Js�a�� Ϸ��<����uK����g�ўº_��\�J3�k���1���h#��K%��r����JM2I^���/����jfr��Xj�[i� ���j�'8����W���zH���-�$&鴍���M����V�ȳW�4�Qg���a ڍ=�ٖ������r�wj�<�����.��t{�vQ���$L�����y��u����Rwu~f��jG��L$��P%��˒Z7ש
Z{��{���/=glM��V��8��~��0�s�o�����>�p0�S�ȡC��+�,� ��l�/��B���
Y�ڴ�&Ov��	�A+'F�xd���֮	*�$޹��������*��{�|��"����ݢ�J�gG^��6_ă�^y>��%�?�����{�xH��k�\���h]�S�[gF�9�C��h�s�Y�.�E3V{��{8��pd�N!���Ώ$��2�/��/RE�LN����K�yE�Q1����Q�A�Kw�,�+�>Pa<L��R�{�ߡ~�`8�fi~�<�4t��W23��n���Z�2N�4�˩�HCl����]��&](]˻�#�2����P�1�Ŕ��00#:O�
Q'��U��A8��>("EjJ@~�hM��<e��@�`�4T:�6G_�XS3�iUn���z3�;F5u��8[��#��6��*��ɽ)��D���R����f��PJ=��ͥ
�s��u�y�P��)��H�,;g��1{f���Lҋ�Xɑ�<Y���P����a�/ȴ�)������l��f��Kj�l>V�JxW5�s��5v/O��VT�����ǲ��*�Zf�C�eOnV?HP��sr ��>��ڴxCy��N�j����#�`R+yĝ�`���v��X���&����ٖKR���ogC<����b�M��O�]CL�֑��<;�(jh���N\<���-*p �����1�@�1����k.K�!�r�D��޻���a���7� �tΑ|TLv�ض;}$k7�lx�e�����/F���Z�?��_��3J��d�^������x�}G͐Y�B+�-ď�x\��>'pY��\�i��͵
3-a{�ͽ2:zXo\g!o�BE��[��"ƴ6db�P��fV�j��Pʲ:�!���F2�o?��W��q�o;I��V��*�+��D�E�&$��v�pZz�u����9���4*,,`~��X�� �0T�a��=̡���PB�d"3A����p��g��Ǐ��7V��Hg�q�d��[�^J�R�
W�#��c�h�o �TMG���.#	���}����y�P�y���z/:V3��Hh�*��h9~C���H\ԟ��z�DS��N�,�w�]��@�W�ц	�X�y�I�v��8M�p���+
b�h7n9�dJ�I�&l���.B�(>o�|��f\�2�����ږ:�c��[���J�B�f�~ӛ�Q�O�\���ޤU�J�T��<���OحiPUx�����mr�6c�(K�"�w:���Wv%׻T멖 �s�$�d�M}kX�}&�㴠��鍊�f0���^ ����u�}3��1�)��T�w�����`M����%.�����?)�1�ȘKm1�l7�+3��6��E�U2�G�,y�����)&�d�5y@���&�Ʉ��.�����Z�s���EV���=
o�Z�<�ƺ�S���x�������\�e�P�-�Όջ�����s�|�s^�&��R��]^cG���q{Xʯ�x�d2Sx�N_5~�]�����q"�B�T:]�z��t4�X=����g��V�u&�,�6���t�X(�`=/@ʨ�ds��%�7��K{�	��=��zpp�1�(�gU���QM��4�A\�"C6%ph��Su�98���^#�R)dg�4���n��9�8���qg.gv/H����<}2j�ٽy�"܅�"e���=�Lm�ܷ�]�,�lkn�hW���b��z�w�匐��I���3�a� |���]G,P��_�e���4��ŵ�C�=�-�����g�'e[o�&�s���gG!�
\�r8�EvSUu&n&��`S�xn`:���K�4p1YG�u�304`]��m�`��CU/����s;`�R�Y3�Ce5c��D�^� ��a�m:�9��?���{�vZߚ>���տ�ԅ���p�nr���X�t����:L���l6��L��ڠ�o��3��x$��{$^A����L����;޾ Mv�Qw�`Mf�����IN VԬV�3�������o,���{;�wm���_p�& �U��Z������
q��:�(�v:V�|�W�s��kN�1�~(�:]�VZ�R[p��F*��
��e��[6{J�k�L��Pg�>1?�=n?�l�2�]���=`?y��٠ʯ5�	��"n�h�0�o�fl�O��M�4hr'����{�BO�SF�Y�2Me$ٸ1p�>l��&0� YR�&i��J!!��4L�R����.á�W�н��O�M˃f���S�_��l�J	�H��N*!'yrpF��ڐ��Ci���B���A��Pyz�6�d���N%�O������6A��δ��Y�tEB�2�0�p�"Nb�=��������\���I�X�/0T�d��Z\�;�Ϩl�0)\Y5 �$C��X�)]�p��1���&]cx�E�?�#y	� ����W��C� �6��w_n�D1CZ X�[4���HP�YNH�K_�S�C+������U�RO[��޴���7r��_tdU���S�j�Q����<3��T�������-�Uw+z�U�����b�X�n��t[�� l%�eHng<���<��u<G���i��0�:�
�п|=ڮ�Yߧ1d��2SmOj�n˸x�Ԕ&XZ�Y�5 w6,5� �ڛ��'��{P���0�p�Ki%�������po݈�m��/)JB��'/�9?X��=��	ѧ�J/:6��U&7PV��+�u��gj�K	 ���>�j�Dě^�L���׸��<Z
�E%74���zq�u.���R~'F�)��q����7�����1 t�{�]	��	���FI�p���)#�Y;y��QX�l�#D4H����������7q���w�vZ2�(�����>)ƾ����?�,>7��s�	�I���zc���mbd�QHD:�����,�v5��x�W��w����sj����0�Pʰ�=���*�{Vkǿ<�D�՚i��7_6��]���B+��64|���8
~;�D�p�Q�p�bK�8� ٘�����f��h�v�������%�]-s��Lʡk���(�ٕ���_�_���jX[��D�Vۢ��+6��\sލ�ڷǩ,)?.*�E������2Ş��|e��F$r��̨F�y,25���D`��pV�X3�6]ְ�C4]�k�c�{;P��8�9��Gk^�u.��b{r�?��S��az��-������0��׸E% &��Ǽ�d�^�����h