��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V����hN=��a���)�硹<H��׮��`̼��D�g�;�mR�#rj��S��k@'�q�/�ha��pc�R�(��g�F�ו�����`d%D��G�qK�DW�+X���iv�O�O����9�t�0���`�<�F�2MGJ�g_Ю3����Na/��4-^}��ru1������>�9��& c�dN���(�lE#�SÆQ�G���-�O�>m�ns'�G�$d�r�S��=�~c{p�Ç�2y{�tڂǨ|8�vf j����o�r�I>�����R啩��E�mp�a��\��Z��#ok:ȼ��'�-%�*S��.杯�W�f���G�D`��t~�7"���N�M���l���ݱ�
���;�a����~u{�s�2������Q�U0�A���+H�L�y���{�Ԋ�x����; ��������j-WQ��
S-:��� ��kXr����7BI8�A��4xt�?RxT�c|�%C��/y��y��%h�f�Yj��������/��4�����T6�.C&�d(�g��bƱ��'�b:�Ψ�OX���p�e=�s����g�8$2���}�U?�C�����>kol[|{Y.ʅъ�#��8ž݉S�<�㍗�G�`;�&���� �P�,��heK���E/L;M�4}����?1�MKё��&��a��5�2�6\$1o�nH���T�LH�ycv:;3�:.>^��H�8��G��X6KԡAqާȲvY���Z�K�@Y��toa��w]C��H�"-�"�X�*�TD�<$s0�-�o-edځ�`���\J<��q_)N�{�b���LQ���|Gzq(U�8j��5-�w�'?����H�������̦�8>�
��t �-�����p�����XJ�������+��H5:�����v4���`uТ,���+�!`�ݚj&�Ǫa�Ĵ�б� �,��g�����b�>�T2�֍]a<o�nh#Ę�o�U��3$;�������?�ˇ>���Tse�u	���$�ݡGn{Z#�F|2g�O��+}$��R8xR����D� ��~��~|�Y�����ƀ��I��A�?��w  ��:n��[�db�Þ��X�Wި��&=?�%n�{,�&F����?��#��-�me��(;D�����
-�#�K�C�$�'��h@r:������@�.�ܧW��฾�t��Y�Z��t�/�h{�T���^��YoLD)�o=�ඊ4k�% k����ߠQ�.����Ȭ���z����1�|#�S�v�6�-,\��S��|���3h~�Ck2���a��5��!�d#M�l祃:�AGy�ꅽ���GD�,yۦ� b�U��N:^�Ff�Z2HGK7����A(�)�J����͟�4�l�%4����B}�	��, �晹3�.و�f�*\�>������ ��K��^-��K�r��\� ����,�Ox�
%�H��sk�&� �K7�.^bI���΃ť�^�2��	q�"����Vi$������= �����Z��j��6��5���m-�"ui,S�ӳ%��m������?��Q�W���12�I���F�Jڹ<n�P�w����/��A�jz}�I�����K,�Q�����o+gB��[#�LR{"��zi�[��ܾ�v��1qc+�J�����@l�����q����������c���-�i}����չCW?p�J���X~�JǸ�r}U6z�?�D[����+���1�]�T�L���{��@�5�E�Ho�w,��+"�Q�C
�( �3��T�cu��T%�����px��)����y�`(�91�[�>'��>�;4�ꀭ�5H���6�D9��È�o�~�9�N����e��>�yrS�J�đf�0sD�A~,k{S�ZdG��	��[��s�A,E�}�k��y������^a�:9�e&tF��"�hwF���W��vP�u���=�fƿs~��4��=�TVmv��=�j�7/_�m=E����PB)sR�_ ��]0/���s$�4�h�z0Y�,�x��Jb��vKPzN8CRn��s�G�����Se�"��}�&�r��~
��Qڅ�f��*1�ه��)��H��ف��f�����p�����V& _���b%pЄm�Ұ��k�ѯ��/�4�
@�V.~�ybXj)�2ӡl�Ӥ���S�x��TyW��BY�y�(��R�mn�G������ ѦU�I�)56^�:"	UB���
�63��[���+����F�Y�E��`׍C�.��B���"�R����G
9tcr�����{xQ�=w{dE�B��P��ŀh�շ*�财^�1/�hQ�������Q�O�p�o=��=V�k��0�↥���������½� IE�S�j��U�v����6���p�R)�C��m�O�&�q3�����u�ف|$+y9B��^Ma�b&�7jtx�����[���m�`�u�F&o�W���'�эL2����Qm�k�Ao�Q���p�Ǟb|�0\R`�
����'�W2��਷p���^��q�_J�� �~v�x�u�x�:�iL��H_O����`��ufVK�����HN�l`*��9;9�W�_��@���B�K�K^ƍ/�^�|���T�組��ے�{��=�C��|e2�f�-v�W���)�G��xd��6(2��]�P�!܀&FuP�j�{�e,b�;�O=:ao@��^�y��Ti��1�L9^	m9�F!>1E�^&��˻�	�qyR�nqDWs�/f#r� ��8����լ��C���b�%�	^z�旂���^EU;��/a;W{F;pr�<�YI{�>a�Ӗ���kBQbl�Ĳ��u7�{����ȕ�fY����^��v�A��k�w���\<��Ь _�FN�5N1�k���b.i.�����f��g�l.޽O�yt�&s1�t�J>� L��~h���MA%�,1��9�z��K`��g�+D�q���o-n��>��g�]�ZO(����(X�"�â6�~���R���?8/����I���E�7a*�v�G��eT��=+�ݾ*HG�� 7�H[<���!7s�B��Ʌ����^�s���\�RK��
�_@�f���ǠCP��m��L%�ɲ�2֮r�/���mL�Mo/�_�2m���[c�>�@/cL03R+?(ɱF�Zx�gl����8,/`{���Z�$ʰy������L��C4�8�sm��Z��nSE[Oxx(^)@�&��+dP�!���H��L��޺�!�Ts��ʙ�R%KX��0\B�m��ӈ�De2�\����� ̆l���*�ıZ��+�=���l���e��U�`�bo0�I3:K%���TcA vإ�ٛ_7y����G���56����gARx���3kI�K �eNT0j�21֏$7	�y���S�]���Ю�Gya�(�Sb-j;�k������!$�Y��Td[��n��՘͜%����~��]��?d'��+���uOMOLz�}˷F�K�F�q�*0+u��̦h-�"N]~��������(�i
 �{��:Q�P�`�g ,8iaY�
_���ԡ�p�*�ְ��@�Y$�gVO`��ҫ�i�Ͼ+�u
`�����@��ͅq�Q��ϡ��b�֯�|y��a��o�l�5��h�Yyղ��Y�	icp;���q����~t) �����n�|�+��П��ֆj��H:y,pY�:�iLE���q7��BQ-R�I�o!hO+k���A�.���V}��<����lM])�����]�����{0� �K��ա���&�