��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V����hN=��a���)�硹<H��׮��`̼��D�g�;�mR�#rj��S��k@'�q�/�ha��pc�R�(��g�F�ו�����`d%D��G�qK�DW�+X���iv�O�O����9�t�0���`�<�F�2MGJ�g_Ю3����Na/��4-^}��ru1������>�9��& c�dN���(�lE#�)�<�$A3*�qy�)[)��y�!Z���v;[��S��g"�@|;w��q�����p��3Fp �G;�Tѣ����N�Y��E�r�E����^�wbI��x���@�{
˯�kdz��dQR��[�W�z�/s�:����;�V��/XT-�Uo]���ж{a�r�g ޼�5�j��@U����_eg�N�%�Բ��U�V�C\!�	�<"�=d /ߡ��;w�ͩ�!�[S���	�������q�i�H��۶�qҸ�O D�Pz&[���?�d�u��߆�x�Q�n��J�� ��˲�{sk����i�D���;6,�_��r���QA�Π3�����D\Ji�c���S5���t��/��Xx�&T�>�9�k�_{�`?�Ku~8 ��|��f���o�[e�
1�8v��@;�	W��"���c��K֜?]�b"�bkhG)�W81��O������uB�8.spy���{�n�\2/��u
�D���Y��|�6��kWQr��kaT::Ͱ�)�	�
 ��VO�aҬ��]i宽�.\�Ly���G�z�$A�,�6��H�g���b���?�Ůx�x=��=ŵ��j����Ypm�$�}D�9�U�p�������.�'
�w
N����C�S̷����mb�f��UQ�1|\�8�Q��T1��{>��~A��'<iU�UY�r�C�)ꖆ���Q���&�/X��9#q_�y��EQ��@����w`�Z6���+����4�͆S����˽fa�(<��"Np�埬�j�mt }گI�s��F�}7��� J�ħpW!�A~5�ƟM�e0q/l@HA�G2�T�2�]�/�1���-��D}'�����DQ��km�=��B��iL�:��儠x�z">�s�����+N:N∷�'��g�Zo�V��2�X	6RB7���ZX,N�t7ۆ�.�9���Vړ�ϟo�e
�if��.�p�pN�Nn��Z�t�1�ЕWL�"`��0�m���X��}�رc��t�mAO��x�
@�A���^˧��[2�8���|���h��6�7R��{�h������5��*�#�*w�$�H5@��Ϝ�oͮw�ڶ"���	nZ'&e�t��ܩ�6�d2a�Z�7�_P���VP�#-*��,�2�r�9p�ox��q�X�F-�k�誹Ej�bq��A�N�v��y'W�����Ϡti����Q��<B�E�Q@k��)���6@X�|IUuW�a5ī��"���+�.]ﻊ��{��>�����0�W�3Y�{�(�{0��?H'􃂥�k ړ�4�. $ִnm!���
{!��������,ۭ�I�E4�֝����M$���te$)��<d�T�h�-qR��9�J79t�d�ߐQC�Q*�k�xuu�UJC-Y�MT4;ڪb:j�%�nh;<�><���2�nS{�2ݷɌ0{�����̃�櫯�tb�����?��TرQ��<Z65o�8,�^��ڽ����͊���3d@��t�т���*d� ��E l_�4��\��&GɞME���i.ZR,3u,�H��[dLxL�濾Yr�O+)�g8g��.��s ���H�
(���2~e�v>�F���Rڈ��k)@�ga~�"?�W�!�;�r�X�U�iW.?�/��D��]M6'!PD������/�ia
9�~���3:�;��_�,�P6�r�d���� VX�ͭ%f��xdv������s{!����	p<j�%�*Dфs����`���������.�#����/,�{�v+;J�,�e"��^�;���HO�\��V;�-^Q�#Fb��0=�d���V3�҃��I��=�Oy7c#ޓ����_��~qw<�N�� ���u�0F��X��xZ���J��͹c�n,�tq���i��h��*����©�����LV,Ρ�*�b�F�,�*��͌M*^Ʋ�+ɃWG>[�Ƨ�9��D�P{WjH2o�<�}x�|���t��)L��0;Ê���-��b���h7K0�r��'N-TFݢ�˪�Bt��5@�$�*_�p9���,<�:�����:�Pކ����*��	#�1{+(P(������������*/r>�f�����6ّ�v~�Cc��x�Π>��*a�$0�J?u�+���G��[W�I_��U'1�Ih:`���D�>�f|�w��
�*,O�5�{�	�v]4?�g�7Y��Rwll���O��Q1�
`W�P��L����mJ��g�����T�q6u��������WQD���f+��^�����f�%��Ѕ��� '��A%k�&`�`o����9��P��oT6�[�-
N�J%[���#p�#����t�
�#�����W�y�
iz�os�Uό��C�6D��E��5�*~�)5�*�u����"��XS�H�]2Ȓ�BvbN=�=�k�Y���� `���\=��HT �3�v�Pqm���7�A���Shf�����h��ht&����ԩo��1M�o���g��4F:��d͞���?���2*T4Fy��saQ6��L��z8������~֛SPO�_A_ߓ�r ������\	-svL�y{�D� �åe?��w��B-kON��
KDպ6�y�I�s�v�K��ɿ3� ��l�]#v�0�����|�}`�o�����#g�}��nD[cS�_�&�q+�٬��dG�0A �e(���>����m�&<�b�N��$���J�ˊ7t~բxc�&��������mhI��V�SF�7]h�*c�H��,��*ouӼ�D�1#3��'6w��Ⲵ\�K��Kb�&;a�R�?�<Ȓ��ű�+'z�a��@]�^ckQ�b.� �h�+��oA1THC��yl��WY� P豬���(yK���$Lk9-0z�����~fm�s��yqe�r��>�Ƽ��T׃����ʱ��wD�'k]��er�zHF
��2���:�<��Q
��;���_ئ�Ʋ|
Ĕ��<U]4�S��LW�`e��&�z�H��k���%c���'�p�*Ŕ�f�
ޱz���&)�zL�>�Z�-6�&@x��"`]���M_DD����WSA.w�����K�tu[��U
Ū��.1@�s�yU�䇓� gg��wB����W+���L�{;�Q�CN��4Ԥj�ܹ���4bʲ�֎ .)G>�=���Y"���Le����Xߑ��}H�� !��j]�w`��l`7s+�-
b`�s���;�n�k;��vI��xלv����bb���ǷR
Rj#�ǝ��kXjQ!o�ꃵT5�{G~_]-�b�� �lrI���z~�B�z�b2���#)���P��
�`X����?�r�.�	fM�6�b�SAb%��qh������皝����Q�94��	��_�a��2�8��+pl��ZƤׂ�@@a'`�$����b�	G����}�:s��]P�+��0C%����?9wDO� b_�Ob�IOW����D�lV�3쩸�l��5N'F�W���tFRs�5�KEBR�ъ��Qr��S�:)0����|~B��<�<����m#-P����Up�K��Ԥǽ�}�oŴ�p߶��so��&Ϸ�g�VO�7 ��������:o��M�����eĚ���?3��1:*����揀�A&�\�E���C-���w�9�S!w{��CN��/a����~�u\B:�y݌r!�b",H��vU�x}���U"f�2�8.P�8�&���
^[rM��9� �D�P��g��.�Yu[�9������STo<C�K��LH^�&c�����S2,�$�W�5�/����njC�9���wD�[��#9��	ݽ�OG��bE����6���q�8� �}�P�;�	���-�� b�q́]+KS��'�)U�5&��$�al�}���z�y�l�奸*��l��r���D�;�8���j��N1H���G�s��ՙV�����8<���{��m�����^�״|%�4�E{����8Zc�A�0� ��Z�V��#9S�i���nh0�n'�w��'�ۃ�n�G�M��ߕ���Y����[U!Xy��G��Ł֔��ECo|�V�0�1w����y��U�w�c�΂��7v�؉�Ehu�wn/��z�vx�b,��a%�er]1�ʆ���q��a��#��O�&'��[�=!��/X\9�0986�B C]�C�-���Y��Gc}��+�����hk9I��1��C��t��U���h�a�W5�N�Dò+@���* �Li�*�P�G��i����8�Ua�X>^�1�9��	��HO�X~�pַڇDvc��~7~����X����F����,xIjLllQ�N;
�sσ��dE�c��^g��'{�a��[�jh�6�P�q�M��ɖj6�(Y�~�J�(,I�V��3t���w�)qW`T^yK;�T	x*��V�;��E#i��$��V㽷'�*�'e�*,Dԥ�-��`�J�����vp���;���ZOWzr_!�+Ԩ߭[J��-ujpMI�,���L��ғ���q\`�
��K�࠲$�aEG�H��/�j �H&�+vEa'���7�EmU�E����=�##I�"
ltR�,�;"ͺ�����d�v*Ꞻ�QFm�䢇C�H��ep��1
��ɾ��(Kf�N�,� ��hjPC�/��ՠ�����<P�Y8�SU]%fL��R�GH�W�I���P/u�A�˅���5�Fb�h�U_��X�/�F��'��]�I݊pIG�F%�S�mJt0$�L�+,�<��[���՗�1,zsS��H�e�ޙyA�EL+eR��z{�i?���"��|ƟN�D��%=[�ukL�V[_"�^=SR��=��E�_�غn?j0��HZ#��+>�jȃ��~�G�빿�ك�uӆW^����	����K���|���גr����ҩǖ��!!��r��/!�����v�R��;�	��LoX��A�ߠ��LXan8�/��.C ~�y�Nʞ��'�/��L���;_�ք�|��u'��Ӑʐ�E��>�L��f}�EvEDf��A�����C0��e/#��7fEf#aW�N|A{]�Q�$��8l��N&�=�E�K����2��u�A�3^� 	���c\��]��i+���a� ���i>C?������ͥ���f{��F����y��Z��I���Ȼ沐v̢�%ni���Q�K��.^"��|�8���.~�⢣8�q���7���͏��'��EtӜLHEX�8��r	�=?��W�F~�����{Hj+��}��!��SI53��7L7l��;J�Jћ(� :�V�u5E�Ʃ΀�v
|�2�Ő�«b�\�;0��ٷy�c�~�@�k��& ��I2�W�c�9�f�JP����2�~7Z�� ���dM˘��:��>V���2��|ܳ�����2k�X�$@���5�WK�I�{p9��os���Ud�ǹ�L�a���rf?�1�X�D�Y-ؑX����[�ʘL�ώVZϔ��s_���I��Tz4h�X�mD4�<{�(�eS����޸�&���T�9_Ӗ6s����Cy���X�[��petl@����D�S=��Ǆh���/���e�7:[ �o C���Ƿ��Q�M��`b�a�6�4�=R�'V�NXHu����a�x���n%k����~�,+6��	�Ӫ�3���o���@�β�WC��������{X�IZ�b?YԊq�B��z�9dF��ޤ�{`�j�/����B�*�k���f�Ȥ�9*�ꎖ@�k�6n�;@�ڎX�h�S��[�8���y�v�A�����2���և�I�D��}���,1]7��Җ�S.�mЦ�O�c�N���E��.L�N��!��c?@$��>s�G��m$����>�:qU���<�.�~��ځ"!Wr8�>�Tmj'�i��5X�Hb�,�����L�c#"�w�����[v� $/oM����� �L��DXr���ǲ�Z��$O�.��o0s��_ƃ������ƽ,��sϭ1wi�N�:,�T�W	s��Ez<_�C�8;�#�8��^6��̽z)�����/ �&zd�ӯ��j��k�~�Ǜ�3��*͑����%��a��� ��Z�PkQ3�:�*�i�])x5h��u�K�����3��'6IF��Ԍv~nK��2��ڑ��ef���qZ�:v��'� �}�	��6vzP��5�F����e��a`F="�Eg� ��z��lh��[�t�sK|Ã;c3��T�NԨ����7������t��ad Ԅ7_4t-/8A�uQ(@�Z�]�*�'��0{̼�2*�4����C�-���!�9��u��l7�-}�H!��*���g��AL3���;��xpNCZ��u��16GIJY����ڬz��N:��N �ʉ:&�Wo2J����t��O`���6l�"�dN��B�{�e��a�u�Q�Q*؛�����'�[i���ZP�M.iAbVc���S-Yڀ�"�A�e��1����}y�\܂%�����mG�|����B�¯6�]E$?�;8����6�U4^��Aj*��k*nh�L0�4�;�+?<6��\R��9i�D%�'�������E��h6�'6������KX�p�[�9��ՉU$9�3���*Y>�eA�ʏǲ��	���{z~���*l�xL/d�p�6j��������ɋ���V�͜��s�{<�����H�g��`i�4�3�
�?6�c-Ƒ�k��J�0|$�)����?O� r6j&�������瀑�P�ؓ*�&��]�i8�٭R�x�S���%	��40a������ٮh��95�]�lx�w��"S@6�����b�ӏ���
�)������qy�X��_$�P
�(�/ w��m�V5���Bꢚ��sH���j:ǖ�2w��AM�D��U�ۥU���]��P6��'��d�Ɔ4�ɰ>����-p9�h�lRc�N�5n����<T��x�Mi�f�P���b���K�1�U�C狔�"3�_����G��N>�TD�����-���d��2�� jiDn׮��TXԠ�e��b;-%��|�_�NR��6@]"� |ϡY%����|s(-���Q��Р!cF_uL��v�ZP�P��ѐ(�b�g� ~�����%eu�L��і�6�pwM�e?�3C�X[��i�y���9�������:���J*�BO�J�Pp��b�� i�#�r�RI(^�s����x]�O䍱R���h�[�c���Kv[{q��J;�p�Ƚ���$�(B�W���@�P!�'��[0�e��Ԕkg�9a�0t3�N�w�F}��_^!Qs""v�w<)��k]�m̔��ߚέZ��{�>~v��el�%)`A-�[X�S�����|_�Y�OJ>/$�t[)W_C�S]rv��ar >Z���Nُ\�!j�-�z��@?���ok
�U0�nZ�'�ȱP��Hz�VzK(j�#R%��x�n��[��?ơ��*f���R�~{�>��~���4X�9�%����71�w ~٦p�^9O�!r��D�G�x�����xь��nh��Z��:�W���)
gf gr]�j[��D����7i�\��AH�E�����A�����,�����c���d�������\wq9|�4J9�"xFr`�h/��s=ZLR��7B?�Q1MYܒ۱��_>@?M#*�Y�~���&�'$�n�+�u���J��LX�탃����6���ߦ̿��eC�+�K3�+���k��u�ɰ���*�H��Ķ���E�:�*9V����P���zoDS;��Q����t-��&�݊��&�2���a�:/��Y^�]� �JJv�~���ex�k��:���a�du�����bq��$(F�@����m�m�㜡�����:Xn���UY����#�p��e�`���ܻ���^)���oC<���P���,R�c;��[H��F�5�f4��6���h'xK7�g!~7�	�&u�i!�Y�\�������3+ib9��fY�:̉W���|�Q:V�l��2�� ܜ�z�^��~�f�jVg-�3
8�Mo����+��@>������"p[�AT#B��;�=�͒�v�jE���Z��H=���T�;F��0]�$�T��x����`�0NM�	��Z?��wG�BX�Y$G]��U<������JG��&j�/j� z�p�8��_�|����&m��@"ɏ�7k+nG�)��C������O�0�L哓4�7���.w�Z}�y�:��d8�(<�2�����]�d���~b��d���4����/��و�C��^�F�}w�,��*��䶯��9 �s�����7�Y��N�e�c)}d�)�}3�����C�郭W�����X��E�}!|vGdM?eL��j�sov�2
z�昲J��!4�G?�^����̄q(�a%�ԕ��r,�<�y��3/2�Cg��	v�f�lsm���=�݉[�4��Kk���Z� ��/�ὺ@T@-ѷ�w�
���]N�!_�pI�~,���G�Z��_�����A}bF��r(f��5�5��
���[�,�i��f�{{޹x)��[�Vt�/��������ouKB������<Bo�S5{�d�1_S��:?߉�����Ph���`�&h����Y���p�<q��>�#�H��2�i˝ԭ~�;���cE���8���5�f�P$c��nѺ8����f��d�I4/9����'�-H�ƚ�G�ՙ�W}����>z���R��L����x�P��&��D��zp憲��f/)o���
6���v�ʃ�G���:c��Bdũ�/��X�&h��zm��Ν9��8gxJ{,XN�H�/�c1�#A�)\�e�;4��d�Q"�^�����H
�zo��e7��%�_vA'L/��H@��tk�\B��
�����������2x�i@Gs�U_DN�м:Z��)�La�� �!
��c��o�Jh>ГU��n�|g�@@q����#��sT;^�Oxv"J�p0��,.I�Yd�i*3=y
�5����.�m�f�fgiف5��{�I���μ=����0�+�Ba����{�M��pVo����eʁm4�Yj`�oRA����c�l��/�I�M�U�҆���Z�j$ݟk�����p��]B;���4G��9&'��lڑ+��F+%�}z�����k���5VR�v�cܸ��h�c�Fk`CHZ�L�}��B��")��d<|r�8ZPlh�~��y��#��Â�B� 畏��ƍ�@����ͿF<��)�Y�yWVJ�Y�O�:! ��S�*SViIC�H���m"������q�R9 �r��_�A�wN[T��utbV����2ϣ��=�$���
�����k��k{G`���7.�����^�jX&�\�gG� 4p��hl�Y�]s�f[�h).\��T�싱�Z�b;S�н"ˉZ�)�aE=��*Pw.��hA
�����佱ϊ������$�����Vq�.$N?��)v���~�ٞgR�1�� ,u���n�Ip�極h��M=l|��ʅ\�&���A� U��!t����p��Ң5� fg�=�ȼj�}��h��� ɣNl9��-�0���,�:s�i���l�hu���ߚ<�R[��X8�I�sS����� ��G����.�%ˆp��̇b������v��8�_Vt��`���Ǫ� ?�q� I40L=��t��)����uM�sZ�7�&��*��=%Q��ۘm�+�9�Ĉ�F"Wzm��kWz7W�/擉 ���ӘUN�O4�
�{>��	�oE9U���@ ��!�^���m3���!H9R�����g��F�'�/M��Q��]�L���{6��.����θ�^Og'���F����@��D����Hј�����[8S^N�{�i �Z������MeG����t���V���QD	$�@�m*F�kc.>u�\K~��>�Ƶ���iPZ�s��L��x�R�1%���!|(���K����8Q��<���0��(��4ۉ����V�$s��ff)��ИV��ȶ<$:������>�0� �w�h�|V4�����O2��ccy�e�,���~�3/���uNeR�J����I���Cs��t��J����I
�7u.��,��+���".:�W�]�<��V%�vDb�y.�_b���L�ܛ�<�w�D��n~��@�,��$ߦo/l4�$�a%w��ȈBS�!���C�#Y�ba��@� -d�X4&vF�n�PZF��}��5�9��^��d����`?���Ua���^��ਛ=�ﹷ�j0���|
����ra��:HM����C%Tea��=��B�֖M<wE��:ϋ�;٧b
�+�b0�'4.ա�[=q(X��!��#�66�G�0h2�c�.)2n����R�����x/'�j���?�ܵ�#M�I�踆:X���R{�<�}=���� �U.quKk��ȂS���g8�1����`���cW��к���ݨ�-[��Ёl?��QP�����G�*��f�AGsߓ�*�)"F�{���J��|e��Z?�i��liV�-h�ԃv���w��t�����WIϞ�i1å� 9t�iiB	���Xٲ�}T�Α=M�ۃ=�-*@�{	���Z
u�����Aq�G�V��[z�[@������c~�Ć*�[	Y`��R�DR�AQ��~�xo�\_�vۉσ��^��.IG|�Rm�Q��iϐ�Wq��4PH�",�7�=z�MH�}ٗ�dn3�X�v?�aN�=�Q~�Xa8٧�����4����naY�2���WH��>$���/�]-�J�|�34��BT>@���n�������f�Î����Y��6��P�A|eG)tO�R�Zأ ��W��i¤S����_�Q:t|Z�}�&��[�)�q���P|�⌐\v�>�ϪA�g�" �`ݼcm@�jyU0-���%���Z�sI^���wə�!Dxl6n�i�\��U��<tO�f��6��GH��.{�c�M9��V�0����uVjH�A�f�i���X���V.����A".��0**�U:���h��D5����Ќ�	@œ��}a�[�'�z��������;E�W�} �b�ϐ���z��W���e��&��8īY� �S�����Jz�o�S����s�����o	����^Q�'�	������yA�	@��sr�hv5��X��A�}�, �,�iäҮ51f4(�{t�*7��J/�B`ѐ-�޻�'�����FL�6��@�(�W+�����H;	�������|~�G}����� A�X,�0�7��	Vw>&l����^�BL�K��h5�{@J��<6Ejb���%'x��s�c�e}� �8<���:�%��L]��p.J�N�aࠤ䏬}�ؗtl绸�`l\��R����|	����ع��a�0O�����7�X~����z�/ nO~"}P���?Q��_$�s�r^>Z*h��b�QmL�>�M���fT��4)���l4�{�D�{����.��uÆPCq��:ha�0���{�4=+Sκr�|H��0�|���t�<w���@݌�����Nl���s����Cp�'��O�����&ޢ���0�y�m*�"e�W���U؅�{>N��.�\�kA�Ĕ)@�h�0|��֬�T՟�08��m}����Tl���+H.FF½h:�����"����:�r���?��J�CGӥ7RY��ꗩs�N�J���gi�[N7 �+^�p-P 	�W�Dt�q}�ZtnJ��WD����|�;Z����ui��.P��k?W`��9��l�oM_���h��a���Mw���h�6�`8��>U� Y��cy���v��1[�#"`3������*	��\�S�d�@7�t91�O��d[`���5��	Q!���zW�v��t�Z�����(���^/d�Ԅ�/���>��\L��)'M��A0;��[%��N3���2�xs�f�'�(�D�af���H�1��	`�����*xq��jH� ��e��.JO�)� ��I@,qPzM(���jiP?7��>��%lry���|��z�{YI
�OWh`�� Ue9�EϦ깉�&;��w�\�M��=w? V�uj��:��������2=� ����"���
��.�Z9%?����rv�}�i�G�ʘIi��>E4	u����û�+3zB0_d�_QW��Yc�����͘��	��p�tO�섿,h��]��)��1�m�$c����ч��3�!yj��O�!8��!@��]�N
s�k���6	�b6/D��e�9lFV~p����1���kE�U�zJ��{:�\��40�k�G���u���)Y��wwx����I(�S�h�2V�ʵ+:"���]�N��6U܀�6��m��a�VV�j�x�����&c�Ǉ]����_F�QE���A�`������������c������"n�!�?�:�����J<�[���;��Y�_��rM�>�Ӯ_1%����@��YM-�xM]��I�L����y>ҴK|�F�}����	ѵ��\�C_oZ����f��h����i�Չ6�+Cv�ط-lŔ��CاY��՞�r���qhG�y$��������9pt·���_���_��*�O�軾[��/ɦW�S�q$7���D�\%H�D�A�T�sSpj��*4?�YزI�0G��L�Ƙ�B��r�f�n}�@�RH1+�N ĴA1��hj)^y|R�%G��J��%�?}��ۋ���o���GP$ؑQl����m���[�N���i���|��]�/�p&D�bWш�>��d��7��F�WF���R�l��Xt�E#��-��@B����(�GN���$;8^���0��)��y�q�e�?6�f�	{�	�p]�^:�e�`
�6�Т��R�L(���Qp�F\�$Yݡm�C��f�;�)�A��d��'�O���J��,4mR$��ة27u�X��q]�����`Cdj��������k�i��U����0SB���C5�Fa��ޢ���m/�C(�o��B"���|6C>1��R`���/mW� >~}KN���xw�.'G�B��ܪ�=y�'������������{����(�;G�����)���~�|�α��awoo�G�:�J�l,���:-H�it��-�ټ��	��Y���u�)�m�j����`�S��J�R�kk���l���lq*��q���W�R!V���V=l�E��n�><�S�(��'�Z�N�q�K�n�E�<B�,����Q�9tv�DΫ��<3N�S���m���Yi�H^zI&R[�S2{Ӎ+6����1;�f��Q�L(ݴ����l�;�j˹.�2����c�fqu�G)��^� ���'2?���Wu���D�t���^C�2}���lv�mU��y��q	�/OްM�c�1�@A-E8M`�YO3 Gvؒ���!���8�c�q5�S�sK�ۜCE}X3E����Ч�G�z�uP9�	eL{�ke�/��?lYXF���Z:*?�ζ.�eb��G"�F�0l#6kї���n���L�}��VD�����P*����S}� �֔�h��ԧ��iv�Ik����ݻ?x\5��˱�5�׶O����S�ĝ���7f '��F���s��{��3+NO�n|*
6+-R-��'*4��y ����L�ttC5�S჊��O�&�aE�@�1�
��yŸ�����cS���b̢����n����[��
B��BK[�A��1��	$��N�(e���H�m����}�i0��dx[��Ɋ�o+/b��J�;�a��H�+��uͅ��yp�<J7�CcѶX�)���xd�u!zu��[��`��BN��0&����?�U����Zd��4=������J�����W��L�L�(w0m?�pbZ0'嚙��`f_��_n!��"
rZ�D�	���\G��J�f	H�˺,�$f��+!}��tu�y��� ��Qs�k[	�J��\���5�Qu���E�vd���=��>�g�>����m���m{����`��>�ջW���
�?��#b���S��4u%ɑ�~��H�=qk;x+�����HȤK��$�y��x�ڸ`�b1uv�������,z�i��Rd��qL� ��R���8FC��������W������0K����|��\U���4���/�r�����g��Jx�5�г�;UM��E���f�L����>�*)��B��< ��P��A*<� f�i[/��u��#eN���e}-zWdt������5���'���.r��Ρ-9����Iϊ��Lpې�/t�L��Aĺվ|d���r�3O�G��cl&a;�FZ@A�����������W��XAvC��>y`�բ9R�h�H��?��B�GTP��-�Ą�۴o����Cu �
c� 'w�P�ĭ�^�d6����o�$8�����-/��Z����'��\EfcVE���4���(6�Wj�miG���}~�����a���{`��v�H}&S�p�`���X ]��"���-{��{W�ר�T�� +ాJ�D������n�]3D܇��vb�&ա�<wIŪ��j�SIØRw���_a��WL�p��`Ye(��ӻ��I���L[�0R%�LmC����I��|F���xeD����ߑp�����=�c4��@v@�`�]DV^�v:^� .�6������k��t1]U�?�3CY��S�0���;������L�&N̌g\x�3�aC,h��z"��yA�T�'@_�9d��~iC�)t.!y��C�*0Rz�������(6�#-�JW�Q��T.ܜ&�b�2��� +���[�����������1����[:�gd���Αߐ�ظd%�
T��2�V����Tε�5ѯ$����v��I�QJi���̸B��v(m̻uQ�l�{	���ŰU�| �(�?Q�K�P\�@����%���(ƁMs��h���!�C�����S�5��,�o�w�*��ʅ���ω�[i�Jl��e<Z������9i��M Q�D�^\TUA{��)�E�}��K��c�4����.�b������橙�h�����x�;���̳�N5<�*	�1�W+��ɔ���WCjTC���{c>����x�IחN��G��p���@D�Ż5� ��MoWI���Ҧ�`IV���-�*��7r&�{e�䓎J_�NlWSZ:.�H��d���f�M���tkvB_��a@
���nEmo�@���2ے��֡� ǉ��˴xmB	�en|¬=B,��a��X�MT�=Ǩ�l�k�
�t�i6FD�<C�Q��.����U��7JJA���i���ʳRV��i�XLǖ�ӷ�����7ҟ�5w:L��t��)�Ix�&$���eJY���s�_����e�O�ե�c&׀#.X6����s##�F>L�G��G�ޅ����C�ż�D#�}-^�8

2���pD5 NZ	�+�<�h�g�L/C�3h*�":׎.!���Hi���ɍ��Q��cf*����.��]���|�mPs���+�^��@�Y��:{�e�ɞ���lB���eq��ī!ё_L{�'�;/a`H�T�a8T���ĥ��#F��@=*��2�|mo�	L��<��s~pz��RLrp#(�Dc܁D8"I�rS��x�LRȽ��h��0cc#��G��U���ax`�&O𦏳����-Bh|c��|��H�=Ȼe�$�h�5r`�4�ո��.h�':QTAfT�#���<��m�(�	��ω.D��J�Gz�����}���7~��әh&��ʜ/qm���6]�i�9���c��m���n��68 S��e?�V�z�3��+U��ҏzo�x�+������.�(?ܑߋ͵�����E��0�Uh��Yij�u^^���hnQ�V�����uB_vžѵ��(f{o*�͔w�vs�{u����LN�vFB>��O��2�B����
Iق�s����;����/�P��:1��S�VP>y����kW\�]����[�H��zt���v��(����B��>����5����U�+�yw|7v���<��`���FEKm���[`��+���u�zϬ|�E��т�^>�B�ڧ����ۣ��[����O�!	��}��6�хC��DS`k	!��y��jq;�Z����+�R�m-(��p���^r�JT,M,;��~LD�44��Za� �{�vB3s��Įn�e����<�te�Ra��dI#:9�O�ܧ�%oD�Ff��V�;���~��[EK'n{��}��h��v���|Rk�\�O��ͥ�vJ���BS�{V%O�9�)�f�k۱�>4��h�i+A��aq8%1$���+b���	���cMKI��!�V �$p�MVa�,��F�p;4v�tV�E�����|�Q�so
�\�9��>��dh3�?�JL��^;� T��c�}/i'z%	���6���\"�lNY�EX�*�` 
Kc�p�-j��yŔ���PXr�Z��3E���PRь��
3k4�B$�4�Բ���(�;�e:+a!�y���P�Pk�P&g�#.gW�ě��pGiڪ}6/@(���Pvƞ�������0�ޜ�� N� �c��n���VK�������/_ʉs����5��i�h�/��W�ۡl~ad��i��V ��h�3PͲ}�i�u�]-��u��K����ؗ�� ��B��Y���&�8FRSm��/%�6h�B(� /�T�8%O�C��]�������8�YuJ�h�&��8��ae����s��;n�Ug����C�4L�P��~�@V���%�H7��:�p��7Ωv��t~*f>�P�Tz .^��m��>��fudFY۴.]�D��N����4Yf�Ų�(�H¦0}FZ���xu0QH+�h'�C����
���ZI�3��%E�����orY�\O?�K!��2��1J"����O|��4�r:�Q�� v1#������+�
D�Rpi�����R��ټ��e�.� =l�2/|�x����wO��k�K��(��冷4a~"��*�k��T]z��_�T0�<S򂡓��TD&8���GW<J�^��y���ᨿ����A�������Ɵ���u�lA+X�\�8l�iՎ����d��O�ꄇL2[Ԇ�����;�9#]x��� v��.$F*ȫe����h&��)��ɷ6�7Ta�ܰ�t����v 2�'����Ayh��Bu�����Hd�6)�1�r�;����E�&����>T�;�`����T�_��ڗ8ӡcdg��stL��i[?8���=w3h�0��͚�^��~`,�rl����x$H��x �,T��7� �3�\m_����L���[wc�����W.�IO(��N��`f�n�f��-4�j7jL=����` ��ڼr�n�{����t�P��@:�;C`{�5�,xLzg�#����L�#(����H�(3��M�OC5xs���/�����s&>P2�4�>}26�^E{t���Z.u���-/�c���|���X����PitO��T��Us�{�VQh6�2��d�g�X�5#9�^Ɠ�gX"��"!(���W����J��0"�XUι�n<0�Ն$��#��s���^��#2��Ͽ"�D�����~�����trC[��iŽ;�Œ���D��� �w�B�.l�!��1�r)���Y�s���lJ �^IaX�Ầg �U�S
�p�\��.�S����3_/@�G|}�o�1��$b�Y�u��әC������_{� �.��^�};�;3���b �9�����uGTEħClhJG�TIK�y�VC$�P�ԏqi"�9��.�	
�q��`{v����P�;�l�(oZ٣ǔh�m���\;��f2��( ��?��z�տg�XJ���J�ԃ�4���}�����1L�S��O�ąB�gr^ٝTZy�-=��'�Cڂ�c
*b�����\&x�p�<�,�*�цQ�z�Y���6����ax�`T�[_��v�q��h�J�;[c�?9*Wv%���ɧ�G��g��[^���Ȍ I�.Dċ�wp�G��CE�	�9�ư��� QIJEmA�fq'���v>^�?z����H�������8d;�M��b}M1}���������d����B�T	����d�p�sI�p��_� ��xG�A�&_M��̽U$�T�cO'Y���,{m	.a�FD�?����\1l?���C�bS�	Q@�n�����j7��O����	�	��t��7ht��y���X����q�wHr�,���f���&H&�s��U�F^�L�iT�����SǦ�u�L������e�`xCQ0~�@�P���Z�{0N���t�6�)y>�DY8�/��x �?��O�1z�RYS��y�������&��s�T�L�b�rF�Ю��9�oq������M{��a�v�o���op��48���,�߉�� s�d��G$L���*�4�aO���Mv~����C^���� "�L�� �\m�T��R�<9��o}���ѱ�*��-��������p��C83\���D[����֛����K�F~o/��LQ�ZmQ�� �i��Me���h�W����3��P�5�<y�h�OA�����"&p���"ԞYAu!2��bK�L0l�2���q<y]���X/�PK��c2�fAx�dr=��(�K,��6�Y;ix�� 58;x
�FbJ�`�E	�� ��x�����C��X�h�'Iu�O����Ug۳;�jțQ��	A)�uzj�D��-����,��e�w{ti���P�!��DA�v����9�ֆw�޿�ߝ?+=y�E����CeAN�=z�~b�����ı��0���n�����r��B�=/
���}�DY�ejUp2�`*���%�o\'�xO��|bR�z�&�-k�Xh�O�4EEC� �_:-���5e��
�DG��zۢ�\ꉊr��W!���w�R��K�.�J,�˔�(���M���HD��n�A���ҟ2r��EB��C�&��l.Ldä'*m Ӫ���6x&�?P�r�<����1~�?mJb}���7����Nߏ�I�)�k���&a�4���M�1z��G��ǥ���I�������9�̓��[��$/k�˙o�BG����z;�VY���
�j�;�M�4���� ���ݼ�q�/��
.l��&}�n+���G$�vu�()z��]���bS���y�*�G��_ �'�R���6
�y��Z��Β�O�}
	_65��dKbk�D�w���C�r{�X�9�㛈4��01(Oǎ���X��F1D�"H��3�U�:��br��Ur}M@���#X!��H���_���&�eĈ�Q���v�+�!t�]�ڢQi��'q=��X����*4�2�g�"o/�r�>"�2KXJ��\ltH,���c��S3Vj�]v1�s˹�~�f3a5��:�(��� ��4}��E�zd�
�G�=�)S��w�R���49����|��q����'�b�� �z�臗L�D<��Ѹ@ۦ�c9.�Zb�.�Ra���ҩ�a�"� �:*:��DC���[/6$�frB�. q�[��T)
'�9y�)�>�x�dLU�?M�h�&�ȗD��#U�i�T��|�G�"��v=�|:�1�T>j�������3�1�d71�V�
�C�woI�<��"+�@�4.��.�i�F�=����f�����_`?�%9�1�[l	W�T*[X�j�2N	�I��<넟N�"#<Y<�)�t���g�f�nM����EqI�PU�d�>"���08!�$���3�{�$�2ޕ$_&���J�:�����������	J�J�O�K�y�Y�zE:s-�3{	E�6<��0�u��ʽ�j-.#�m_\�I�z,�0� �l$�F�x�����#���P���V��DW:9Q�$0�4���J�������;i͕}P%�R�>V�>ӎUV��r'a�;��#@?��=�(
{<H¤��`��ը�ԝA�멷
P�����v��5
�]��B�~�?p�w������u�"�X�&+����V���6.i-��|,I�<�Wl2��b�R���G�}�k���@����`.0��M4��O�Y��L�����|���$v�?�{�`���z߀������7�[��s�S˘*"�B*E��M�j^��D=e*C�#ق�Ci2��Vj�>l|�G�@o���9i88:2 VJV��~1��N�ǚ%�v�Hva{��e&-�9
KBw.ފ���>-������[Nv��ӝ�n��-�p9�~L���Xۢ������;��K�J������gz��WJ��O�\��$-"�p���Zu����@ͣr�ⲫzg����{����o���n��F��GlZ5JO�s�R)p ?h� �G�3���w[$�	���J�A�P�����C�DKv���^�7m=��`(/T�X�|��Ps3�Xc��;�
�flDS��o�fr�:9��;���#�����K���,�fK�l�faL�&�d�K/�A�����Hʌ�v[��,ɯ��g�uQb��k�[(b�:���'l;p��8S���d�A�1Q2t� vR�h����zľå��s���k&��0M%���fUf��\�s�<�p�)��x9�E��%�H�D`!���z��G_�/��i	^�����3��Sv>�Nnɩ���BN�JWS,�#�O
�
����y�]��F�1��=Mp��.^�Ksп�ի���ɋYb^��?,�[V5]i���$�q��GAJJa�]*Յ���$u�<����z¶9���?�*���ԉ��	X��	8�k�~%��gX ��Zq���[��=NhL=��9�[�P�c�5���TBrD|"6����y%l�:��(���F� �H���v�ǲ��l�iNU��iG'���T�}7�k;��o�J��d��3/D&а���g��zhv���0H�vD��k�\�()�&����+�𼓗�B���n�l��֤����5w&~���,�j�ƺa���l�A��Z�5��1c"0��ASez'>ʟ���))�EK$L?�+�����ᥛ �y��""�InX�T)�Ӏ��hr��8��z��ɨ7�wW�Bh<��d������!��j.��أ�	Go
�◹'����'�)�q�y��T�`�x8r��wqGYl�A�^p�����-a!������ȱ���� ��h��
-p�f���@>�Nȭt�,�}C����
�MtI�^x�;E�Ť�I�����g��Cc�e����)�!'n�S���ߣ-�� ��{Lُ�C���,E#�p�����{"L��d�XX�u��\f��tI`ᗬ���
(���Ip���8�j2�VX��G�%N�uu���9��5��=⫅$ZS�&0�Ou �ČA�1�����k�L�=�L䪹D�n���T-�F5���Q�H��\�߳����C9����.�>���`vt$�j���e��EˆH**�I��N��1~���'6�g3!����Z�2����gmpAB�d 8��p�Z����^�w���XEvW�IҒ�2��\HC����Ǧsd#c\�V�yE���r�J��u �$��5U�HL�a�L%��6ݵ�5��>��'�X�tW��m����p&���3��7��2�[E�QH��#�q���U �wľU8��0@8S�ܓ�P�Mp�T��Q��)\�E��JS��켱�u���0)/=�_R�n;bg�������M;������*6f@����g�w�t��̚4С������	X>j]QB����?���
�3���B��<t�V#~)mE�m�ܳ���{��}L|�����Z�u�2X�ȧ,� e����2��g)�qQ�v���b��q�$��W���;���T���*��Ns�z�^��d#_�f4��%���ίU��a��F����k�C���|��V�j"��0��w{Ҏeʧm����>� ʔX�ne��W���7f�@� ��g��q�Ʈ�F��~X��&ԇn�����/����-v�X�\��*�mX$<�-LA^��l+��8�fy
E�6ǳ��®�źY��xh[d)g1��O+o��<�1�^=��>_��Fr�С��c�fNt�e1�[n��kڸ(g�E_�X�'^gJ�V�>������5�*j��?:'��j%	���u���Z�I*eC��jKcE���p����(N�Jx�&l;�׵���}�',��&E��=�+�tԂ��&U_�4w�b+��a�0c����k;U���K��&V���H���4*��cdWD-3�i	X�#|moH?=���R	C�z��#OG(�J�gU����|:Ƌ'?�����Γ��r����;U�a����}�����w�$.�,�^N�����@���=�ixRu�����x�BP���D �8����uC�����ꍰw�Q1Do9�G�<)d찢ؔ!Ge�ok��f��J��j�
L��} �6Y��NPZ.H�pK2Ϝ(!��&���&p�>s4�!s���⣮��W%(+�51�-Xڍ�A�|�w�j��uB_K��!�2�4��%4�	�������tdEڸE�b}f%%$�3	��	�z{��}���z�Gƨ{^=�j$uH�~�#]�\�:����0���h=���@蕅�ɣ�jl��KZ�4������)��^*+�+/��5�9��!��wt�̎RZyc�j��Rk����=]�	$�i�B�j8�zl�7�i[�0H#��pQ<��������N��<�ҁ� =!n\SƸ��M7B"�ȗ%��(-�E���/G���IU`E�=�=�p�Y�#0����d)��&]�8D6�Vk�H�jb��[��GHX�ۤ2W�Nf
��182�aX�R��8�89��������
W0��?�Ќ��*�l�[�b n3��0����i�b%�[�dxf��~o��t����{�%���P�NK�{��FKz�N$9�0��`��#���Q�p� ږ���ݦ�fp;F��&���.<��c��U���O���.�|�B v�Óp�C؟rKe�8�l��ͣ@��m��(n�Y��_mHu�ug3J�ֵŝ��v�3�<9��(�5Nw�>캍Q��gGQ�3��y/����Fz+3�m��oJ�O�a����F��	H;_v�`�w}��r�g ��v�a�;����j�3e$�y�T����d�Q�5��+��.ʸEڝ