��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V��wg��+��1�0��"װ��_�����/$j\�4�eWL}�:�Ԕ��P���	Ȉ�P.#�/;�b����j;li��(�(�^n� ��q&�w����+�a���\��J ?#�r�xtܩ��3�}F(P��G�2�H�r5�$�2FQK��@���I\�������ސ͇�,�-�'"U��b�'�(	�s����C-dO#[H��.�N��|�9�>���sĐn��K�A��?N�������Y�j��3�0�!��߽�p�a�7��D�a��Q*c�B�(Ӣ�K҈�7��wB[�U������Gz���\\I�Fܩl�0R�T��-c�
�A+�K��j��FD�E�82ǣ��}�a��IM����lZH�am���׹�D룺�Q�9�6�g�(�p/}J���y�eV�u���\1<˛ʤB�+[v\a��t�_�Wե��g^cu�����R0D�R۽���6�D0R#4`�����_���8�٤(ߟe@�b��K��o~�t*�0H���7�ġ��9-D�e����3#�'��?�����'9a�'<����R8t6�U�}�:{�s�� ��p�[�n@�(^���s��|hr�&�kv�Jv�h#
+u� �d�>\�
U#�H�c�3c/�����^c��kO���􋁹�O=��6fw9���X�ˀ���3F����尗Ư�]\�$7�K��$WR����'�8D`t-�C�*)C� <��x̫,��_�
�9��Шq��qA�
R�eOB#�U�e?�Oҹ)�U�i)��#�Ʊ���K�6�Mr�4�>����5�#D��?��Z	P5�W�8��u��L��#��.&�u�(L@K�L����zο>f8�cq���W������n�{�X��;�Kv=�"��di;�n+�Ѕ�5d�F�I���,�iB-�|��[�\��C��1�R�ܴ�Y1%��RNdN�`�4`}^X1�k�W��H�e��!��}ɏ/.�ٳ�
|�$���A���ȇ���ޖt����a�;���+��2��x��Ֆ|���3t�C9���RC�D����Ki�%͐��j�}��������.T�f��D���R9tX�圌u����9:؍M���l�V���ᨧ2���� B�%�� (�&�U��(��s�支wPGiJ1���6T��;��'�+�g�o�<+Ys� ��\m��?����қ�h�&D#�yT��W^� r��(M!�x�RI�@����"�. 6AB�yc>����<`{ ��,�n��d�Xx�F����$d9S�Xc�o5��o��"av����f��2�����|`��؏<c����9[��q"`��z�H�� �$�/�R�+�ӗI�_���`�$��!Ƚ��"��}��2,`I�w��9�#}���F�#�az�]$P5̕PxZѿl�����SQn~���#ш�)���'���j1���v�aǤG�T){�E�G1�'o]�������}�U!���% �GX����_���Z?I���k`�^=9!�! ����:V����|�̬�ef+_�q";⿻@�Ě �p��M�/;�N��v3:\AcB8,8���q��C����9�����rm�����ak���A�#B�}a67z"��u�}R/��2k�7���(٥�P}�[�ޣ�ݫ��{ ��M�<k�`���!��θR��|CUU���T�5/��e $�!���Y�Nm��Cs���j�'"��%����n�*����A�O��#uXg�\��m�cI�
Y�F�P����i9;��?ڸ�n.Zֿ�}�+���K�%�ΰ�&�M���U�b�вW�߶M�gޣ�2k��t����s �k/�N��r��|a��L�P��KPU3���7�G?�{<Y �&�;	��g�����Ql���}fuX ߳��YG~����7y�$�B�鳸�:�g�< �C1Z\qPQ���Q��] Tnm�\.j��5�V�ZKS�c2]?���Q
δ��8�A-J>R~թQ��R��m���Dr��z���7����ix�	��V\���B4Y�i��� Sj(��+���Bk%�2��>���W�������=�eyQZr��/�ػY��ng��d�����d)�G�w���DXt�޷�J�N������uqCA2h6��a1�#�;G_8��7*J;/���W�#+��t��w��dNߜc�B����{��o�i��`���>Iˁ�q�W<�y��g[��ϴ���~�SZ|l%�|��P;d6���f�a�~�����{�}!�Uv7F��v����ni�O�NF����C�|�wD�\/-)�+ֳ_���I �s�'���1���{F������u7T��"��5/�7"v;1(� �k��	U,l�r(���ސ�i��O\"�S"����u����/�a�'���쎄�xg)�Ur����d�?���쫹�Q�q��C���AW�p׮n#��,�:�8�[��s �����Z�!�*xh��1EaRP��F�`4:�享�,\�ojC��۩ނ�����{�yM��_�k���������A�C����$gVN��9g*j� � �i�	�aC^��_F!�ڍT�#�bK�d_r�̈&K��GC���_5��P5�a��,��ҋ��]ĪX�p�BLዛ62��	�R�J�`�*L[Ї�m�\�����W��Pv-G�~��^zg�R�.Ɲ��n��'��h��ؕsm��$>.�֟Rا���e��P���?�]MmR*�,v�#8�,H��o6R���u��8Mx��2qކG��¤0����{P!\�t`)J����W�!�ʀn���������5��q3
�#����ux�M	݋�Xf�u�+��T�z�è�_�H��ƏW�("�D]�͍ܳ�Ma^������U��|�6-�q�
���ad�����D�INßn`����O��Ǝ��H�O���=Wnnt��\m�䄡���=��01�`��P�%�1u����L�Qam�m�KœpjU�=s�����C�{$#�ۯ���:��y��5�� z�^��5'H�r\NRm�!.5�؅������Y7��Iܭ��I�5՞T����?���MhHÍ�fd烬��@Z��B��{�F�}�ƭX�QyyPo�*�� �E����7A/  �Q�಍a���O�\���s/_�=��6�{���R����8�(�K��B� W��*�3���e�X\;��I��>�ܩ���rS5��{t�J�H
��%�d}]����(6��ا\�7��y����~�1JP�-��	0��u4��/V3�R�6�k�s6�,����<�\0?���5����q�������r��<;<j���ԌG",�7� :@�X\�dK�`��Op�#;�L���w��
cZ����ɕX��T��zS*K�2���)�E	��IoI��_6a�����J�Wz�0�$�
2�� H	������,rܑn��F�JM���&��g&(-i�����6Zl�:ZT��{��⎊x/�r���t �[]|N��)�8C��҅g����ux$�v���f�����ס��A����Kh���7B�Y�8:���A1�����ڍD�(7�	��+1'��[NK&�<R�CnX�sLp`#>���Cj�B������`kf�lA����o����֬,�2J��ٓO)��2Amj��^S�{�I����	`r�w��Pnn��g��RQ����q.� yH*2���Vk�0��GJ�9j蝨D�PBr�rߔ�.�U�?�p�,;[P��S��V�ǥ���dz��F������2p�y ��i.�����KgPd�|v�AsjBȔ��X�~�n+���� � �-��Sxٟ����M1�Ap��o�Y���N�ɼi�x��H?��(�.��e�r��������=]
�a�k��3��g��y5?q�.�e;C�� K	�����F��6�`溼)��=R�aq���T�����R��K(O�c�k�� o�1���}�t��,�D�YyD駫� �� d��M:��L�����u3�;����H�yu���D�v}^sƵ�}�����%��{"K��,H�{�74bL%��
����uܳ��Iڕc7�I��6u!�r͑џ�um2�HWf�錩�gc&Su}��i��ʩ��~��Cк�%T��ieOj0U*p,�N�\��ԔF�q���5�-�����и\G@O���]��X�
$�?�O��b"�����z�k@� J��l����sxȉ�)�������Ș\��v��z��X����O�7��������2��f|Zϗ��2��c.���|�(���e�%�I���AQ�)X�kRO�*Xz�*IoQh\��$GcQ�z��X�t���Y*z��f�b�v�@%ߪfh�*9�(e5��K�_3���k7���jy�$Ns�f������s)ڔ�}]�5b��j~I�D����'�<��<�#d���|����a�,����a�u��:9��^����چ��/I��ޛ���^�h���E���f�J�[��f���#+�?=-;���}������h�bs�v�G=�(P=�,B�*��3Ex_�U�#,�����H���9�[IW�-�9����M��7%�'|�F}3�ٿț	�/6��9B/�,�ToO�[�0�����l7[�N����������I�`����[c��K��q��
Z]���ٜ����ޛ̶-X�7�NE8� �.}]�Z"��:���Es\�6.�a��[��b��3{9��OP�bG�/9��GN=:��uH�F�E��نwK�o�q�y�+n���qcv��B�ض/*��%�F� �K9�[��J�]��$���(K��<�e��|�,��C��P�� ����9�ķ�-��5J��]+>7f�r݀���J�5�����J.[�J����q�qX�����e	j0���P+�"q��C%G�f�^�	��|�����������߿eb����y�M�$��}��Ǵ������"yS$��OͼT`m�V���B�OFIo����V�hU%�����E*��IUK��BA�K��_��>�?���_������?ښֻH\6��0&�db:칥�55����g�7�8�x���<�H�7�Y�ơ.#�ǀ�/C������L���7<��c�����hG�b"!�g�7~)�-z�n�LO>��Jn�f��ڦi1A���[u99�"
N�����E2{̯���4�ٱ�"#1�M�ku�Un��2F��h�PЙݱ�[��H{�j+B��ޮ������͉�_��}'�9��~�rf�=q��1���Z��9� �=��ok�HN�����pHz�x�L�Ȧe�}Ʌ�W�>L%��&D��P@`E��)��'�'2b�e�b��w� j7���T�������
4I.���[��:�MϮs7�%��G�SO��~��N�y\��(�_�$������&m���(�o�iKX�d����P?����J:��>��Z{JOxPT����oޢ�."��v��Z��vIV�e*�ɮp�����t`�Vnr�t�f�X�J��4sR�#���!_B��b�$���f�;BB!�@,.İ2kLU>1��6X��hE�Lйv�����uJT �����<LL�ҷ��Ɉ���f�ז(MXn���Ʊ�f�Z��A����e!��A��ڭif�s�XL�vy<����Сb�X�UA��Tp�.5�`��WT$�5��;��]7����T3���v���岛���0 ��+A�ixA��3U3ey��T)�c�}��4��mu�J���R��?6�{��CŸ*�������������vr�W˔�t{N�������薎a�JU�v���쐇���E_g��6w�QM�4r$S�5#�ͥ����~�C)�)�Us�`�)�(�����~{�cVaN���)��A�pW��<���
�d�ZY<�N6�^����}��E��E2�
26��0�j�5¶�-��₉=���t��cY�;����T �u��#�Ǚ�hGC���"ޛ�tȪ�d:��AG�1�����t]�,#ϾY<��#��fd\t���5"p��E��V�w���@#fRkY��9�����_�A\#�}3�`lm�c幭!ߦ��=�
}�f�Lp�P�z��� ���fg�jʙ�.�i�N�<��LT=��'BJ"GH��Sy�&������HO�������Xh� 0�'26��1��k}ӵَe�[G�wÞV�KD ��(&VshMN�*q �_=A(�����Xڋ�SQ��D#���`��^i�zH��k�Ίh79��c�-�l��móc��z��ּ�{Uo:��5�E�ޘ!ȸ1ª ?�'x�f׊n���f�X��tW�wӀS���DeQ�k-I�۔%&��[�0���}l�=]�f]�L�
�0B0\~�n.U��7�Pd�z(Ԍ8�ɭ��'9�g�=v��kFN�_f*}�:��f��+�KI�1ۨ)@u�"���3oN�	S�ءujQ�]lʚ�[�.]����ٺjL\��,��z���g��M�I�,�'��	�i;�a_���y��`��5�w#����+��=�L˨&��қo����X_�Ǡ� �3(b�Ơ�+!y�7�t�4^��r��{(���[�V{}� O�I%���9��@�T&���jlt�jK�H�W�/���9��7�+³D)G����HV��廣�6߲Ʉ�EaY*�G�.+STf�
����cFM�IR7���D繇� �-�-̧�uK~��.�F�����	����D赾3��`}��E���m�fN�P�R��O��1]=^�����8��B�Z7jE��������G4�+?F&s����q{���hH����[����Z��oTT̜0�� z4���m'R_'G�d�}�c��5���u�k�����\� �}��]�J�
����/m�ќ|MBxb�M�������-���M�Uy��z�Ѥ�P�q��	o��@��+@�7pOكg(=�I�(��l@���|)N�Z��zӛ�V�P\�E���6��瞔�EO��7�L%J�- (j��Fƅ:�'�֘�H ��n�θ�OB���:y|�DQ��o):>�^[