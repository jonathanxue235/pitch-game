��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V��wg��+��1�0��"װ��_�����/$j\�4�eWL}�:�Ԕ��P���	Ȉ�P.#�/;�b����j;li��(�(�^n� ��q&�w����+�a���\��J ?#�r�xtܩ��3�}F(P��G�2�H�r5�$�2FQK��@���I\�������ސ͇�,�-�'"U��b�'�(	�s����C-dO#[H��.�N��|�9�>���sĐn��K�A��?N�������Y�j��3�0�!��߽�p�a�7��D�a��Q*c�B�(Ӣ�K҈�7��wB[�U������Gz���\\I�Fܩl�0R�T��-c�
�A+�K��j��FD�E�82ǣ��}�a��IM����lZH�am���׹�D룺�Q�9�6�g�(�p/}J���y�eV�u���\1<˛ʤB�+[v\a��t�_�Wե��g^cu�����R0D�R۽���6�D0R#4`�����_���8�٤(ߟe@�b��K��o~�t*�0H���7�ġ��9-D�e����3#�'��?�����'9a�'<����R8t6�U�}�:{�s�� ��p�[�n@�(^���s��|hr�&�kv�Jv�h#
+u� �d�>\�
U#�H�c�3c/�����^c��kO���􋁹�O=��6fw9���X�ˀ���3F����尗Ư�]\�$7�K��$WR����'�8D`t-�C�*)C� <��x̫,��_�
�9��Шq��qA�
R�e؅�Dm��h��9e.�#���)� ��?g�ok
���I��{�Ď9�
z	�5j|g�OA����HF�Vu��~�$/���p1��$u��"�ib=.^K3��7�a-�n������y�.W$5�'*�f�o����\=���8����q�:@i�<���p.�,p�� �{�q4Xa���]���ޕh|�S��+8�(�n�G�q��?���<1�K�O��%ͽ��w�6I%��AUu&m����܂dQ;[.�#{x�I{<���6�J� ��1-j�9��>�,�~�Զ�Ż�AJ� I��IW]�/xAʽGmn�J}HF;��e��_4�5�˖��� �����u�^Qʆ8��1�k��ħ�p�g`�z�4bC�+z�
E,�<6��֐E} XM,a{�՚�󕧰�*�s��A�K)WŶH���F�}i%�	�u�#�aG�w�8���/8�n���O�6C�sh�*C��Ǩ�a4�d(�cg�l9�3>��Q��g�C �U��ȡ���2gbo��ѝ�����-�V����R���]���� U��2����@���=as��/��>r�qa��0asJ���w��)�+^�S#�X70"���Vqz��]����p��of����|EQR�3�A�I�4�_>���Q�K�b������K0��?D���ɝx�h7�������A1�3�:���Z��}-ĥ2�C��R�M%24L�pY֧u>{N֘4q_�\ذ��av��y������Eop ���oe��r��>2�bN{渨:�mg2U�%�+�Mw����U��TE��v �h����rO$�^�k���!���nQr�b'@5�t�����V��Zϫ|ޛ>��{Ź�M�2q!�ց�&��^�ŉ �x�	�&h"@e���=~Z�����yM�y�
y"LP˩�V@�R1qj3�)T��9<�ɫ���;z�`~�����h%�ݚ�I�/si�2�q���,-\�! ��l��?�D�xc, ԩ�Q�I�Bј��bs?�_�0I�S�=x�=h KrL�4a0۝�\�ҭ>),k��z��w��xF^��:�pnn]�p�.x��ɨy?�c�l�L��]��J�m�I+�Ŝ�2���k,���O%)"G`7�v,��ډE��5���@͂���6�v��23�!�]ъ�LЙ]���D���|��8{j�%�O�q�b�դ����;�:�h��L�������U<'��ק1&mR-mb�)��_= ]P��tE�g�a@�����,u�	%��Ev��+�Բ�G��W�n����U�%Ep:��H�$��`�?
�>�u�-�t�<��:����O=�����sE�h��c߰��FO�ӯ�_�a�i��H���a?7�u7��#U�����1���8(A�J���#���s�D�1k�o�ֈ���?���_�	и	��UE��E�&~1�Ųo9�0)��?�hkz$��l�x�c�Е��
b�v � ��D�n�<
ԪĮ^�� �h��*h
���N�a�Z#3�A1��������C��������}��S�x
��]�|���(��K�Zo��(�Js���ii�e
�d�D�sU˙Tt�zS��	sK�e��?@):��^ِ�0	9�v^lP�����ty�ܲn��M	�/Y��@��W]+�g�+A�ґO�PF<6�ͣ�؂w} �.7Do��h]�H�J��I�#M]�<*��4��m7�J�׉p��l��ݚ���޴:������;�� 9Q�ꂤ�M�=�x�Z_�q����x����{�����&�@ӧ	�6��T��i���M��O�Z�xK����G�~����ϒ�������fۢ7qYfiT����Kn�%��3+�N��9No�N�C�Wm��}��c5�EHu�oCH��2�H��"q��b6�W��F�������J9u$�ed��(s6��Mi��V۱
X)~��B� 6�$ĭMĆS�\O��<G��:��|�IV�_t����������l��Z̃���=����?�b�������|���5�I�Ĕ�S�CO��N/+�߬��l#|d�P0��^�P(sJ���A�f`6zaM+")��~��*��$_ ,���$^~���?9���ݰU/#S�����e���m���{]�\�D�cgH.Jjʿ�5`sa/�bÒC�f#<��i��5<�� �j�3-x���1���C���k��g �%j	��ߴ�@t[K-�#Z�����ȶ�8��[�>m�NܣXB4�0mށfT���}��N!(7�o��'\��Y�,+<i����3�����&�Zr�d}���+ʵ��̹��˴
C�2"*�ɭqIN{����Z[�:�J`;�p� �F*m7ݴ���;��.�L�\�ߪz��\k-����L�H�}j�U[O��C;˥��7W�Sv�=�_�y=TvG�7ÊÏ��T6����Fj�55��Z��Up F��.EU+��=f�ˁ� �䮍6�0���[Os���u�rs4����h|��QW��U�\�Ӏ�H�׾�.�D{��X#���8־C�L5)ځ�B�K%dW���ݿK��(��R�`����uѮt71y��U��ѳ�&�#Ҿ%ƀ�E�<҅�/rdP��pE�<�<��sq�5>�Ic���K��L2e�"��N��z����k�&#i7'x���{�?,��]7t����dE������r���'t.���t�O���Oɔ�\���Z��*��_�zcӱ�:���T���`L��W*�[��lL�u�6����8�#��@�д�$�'1�4��E`���W�㶜���M�p����SUbB_K���ې�$�d��u��&�(vÁ��t��4�oƑ �ڰ��')���5��x�7�!�-58�E�~x�k[�X��c ) �~?qEX G3�F��(TװgU�U�}����K����D'}.V΂�_>�A�.�+$��P��1�����)?���E����\Ƌ�w��ŵ����u�sH��y��]�
^7��ǻ&eG���D�Kt��DP������s׍���eT�$�������|�e�����	�ɽo���̃���;%S���A{#�"����_qxzv[`t
[�]9�� 3b pcVS%ˌ��:�������d�!`м��Ȧ���dS�?����9\��PO��� <'ţ1��`tA��B��C�;���S+�y=X���v�Wt�n����f�b��Vw����N�a�@���j�Qt�A��\��
���Q3 �:�]f�g�dџ�v����(V�|N!y_gI=bC���Ε���q\~V��>x��0Տ_Ő�$X\C�C�)���ܟ >�RQ���a�S������Y�~��{��V��~�ykI�X~~M;���Fg�z�(Md\x5xP�����\R�JO8�ξ�d�i�s���C��h�o�̙\��C��C����->�]����Z�S���(�t�F\� W9�'pN�$\J9l;\\"����\M6� ��4k9f����}�2�6*��^��;�9c�v=����5	X����PRbZ~��j����X�Wu�x�U��-B0Ba�|uǂ$�~�O{�\�7��i��Y%���G攑�|����KE�_Lb�Y�W��}�3|8[�@��-�_�BW�i%����(�+"MX�wx������N�$*L�~F	ddU��b_�S�K<�B`�Id����%&�;$>jX����%�]����Q1J��������r�g���� 3T����蚼�l^�^���ϻ��E�>�ɔk�ͮ��w���ae[��6+�ozŔǛ�}�0F�A���Ɏ[v���Q���p�XW��%&ې���l�f����F�Y��Wr4�@���% v7��&�s�#���[%1s
�XP�=�_S��a�$=�X��Bgb�U�y jS������`�!U�;��U���Ϡ�OatR�����Q���q�x=�e��OA�ıiyD�0�U,Z!�����L\2��x��W�,����M :�	��h��w�j>��-'��n�
f���O�/��^´* Lfѻ�N�ߧG"7��*�xp��G
���M
�����{�A��u��I���_�8�NR�;$��G�=|����yj"�����ԫ7�@����+<��w	�C������e��N��B�o3P�B�(���܆���C��ab�e�š1#-F��Ly7����~r=snI`�A\�ioA�
ڵ�lu�ѯ;���!�b��Ĩ���j�?P��m#QcCCI_P�&���츇��2o��{k��bX���RF�#�ʌ;vhq0I;?���j�a��pY�kp����Vp|�S�X�A'g+��$�ȱֲ�ز�v�j��R,wn������3�9*!�ғ��0b{#�+\����4t؟p?8p�a�k`�'0)�=�\
�:op�{<����̨��6�(��_�R�q��2˄~DS�%�}Y����h����^	p�8$�*��[��yp����d���b/�>��[F�Ub-�+��EDK1*��g��ef�~*���@X�Gk�d7��B|T�������쁚A�Np}{G�]s���7�8[�&� ��-҇p7�Y�0hd�g��E��~�!eT���'1�!H"s�0d^�~T�ݻm���GZB��k٧���( ���^[����o�����f�aw�OU��l5�&ek�piM:<;ڼ&�6c	�u�S�#ZDU����/u
F�n��t�$1)�T$1���P�����7B�0��{W`1��[��f�QK����!��e�z<��UȦj��iMt��;������9}����
	������~�|߆�l=�
c6��o���0;���`^O�&TÃ))�D�s4n��$i�i+U���:��70(����.J��B�%���M-��d�lw�FղO�{��D��^6��zb��?$h�z�d��9�����CUڞw'e&�c���nks`�w�_t��47�`�Ҽ[?��7ޢ��2��]����8���b��K*�W����'�	���l8��1��S_gՂp�$/�Ҝ��I��m�$2
���.��0�
�t~���G�|�ׁˋ��b�*<Q�a��������Ns�XW�-��J28��L���V�m����q�(!9��s�;�B�a$m`�>����&�&ƋK?=]��q�����*�hZN�[�Z=WaBywq��䮋F}
��u�ȅ>���^�K�r��WJ�tw��n^7�!+���0y�X�N~��.��*��D����-I�i�[���xFY�����嵤�
�7�ϭ�_Զ\1ǦA��cxM��^�(a���}���	�<Op�`� k7ٕ6C��Q,��@?ܭ�W}�SΙ������n������Y���3"������� 	���cRV�9_��z��~�ob�2�g[��x�J؈a8րN=��+? ���&� S��ݤ�
�+�p^�ENl�L��9ܶSp�'�j2uB 7<-���l&��!k��b�)�^�uRƦk�0EJƈ~r3�r9q�Ƿ��k�b�?&��6��D��4u��4k��9ļ�{H2N�;��-��ᗄ���������t���izƏ �?���{�jVCl��M윗�o�u�M�������}[|&�[����]��Ac�,�Y��g YFμ�~��S8����MK�D�y�wVf�S<TD��9"`LE����<���0�8��0:ŖZ�WhUJ&����r[���&�.ӝDҎO;�Q|��"��Y�����{#D@���-�YC�(r�d�qM{� / ����'ߥ��B(��mӔ�H�LF�>?v[kX"aQԪ��Zό����KiL�|FK��XSW�Sj��[ש9�]������)��W��
�V4•T��5�i���w%Eϟٶ���E�@'�����o�h�ë��[���ˤŗ��fh�Ǩ�Z�sō��-i<�������_w*�H4N���މ������b��\���fMh4U:Ѳr!���3�YDI�ѣZl �dI��u���K�dəH��G�YEW�[/�;h�M󩛡�p�v{���ݠ���Y䎟%"�ɛfi/�^vG\7X���R��ɧD0)�ET@�0^:�a��&͈m��L���C�m�����/L����.��J���!�����	����#�%�"��;�W�J ��7��O�+�w�j�U]{B�G�-y�!}��cW�2��fl3��r�p@%w�����P�Ͼ�0�>SgB��Y�a��,�ԭ��E���J%��}t>��SȠ�RV��5!�>F���␜q�[zE��� �R#e�������r��p�A�{�r[�p���Ѳ�}�k��櫤�?Z��J��w�1��V8�;���ZX���X�� ޚ,f�_E��:�A�X�P!�����a��q�z�O�\y��P�7EQ����p�O�w�x�k/I��|@/����>J�ꂂ�2����J�h�]�l�'Y��awj}�X���r^� E��$h��Y�1�OB�?�^�l�?����Ak�֙�$��b�=`�g�S�:��Xf4%��Je�$���/�X�-n�6�l�� �(��>W���:����0�_�P6%��|��%�����C��sU!ג�_�������n8�sv���!��
Y"[�H�G�����#�/g���~`�zV�Y�楷�/<�E��c7��Om��@�]���t\ (�7��(��VB�l�7_V��v�����ī��@�<���q�#�(c��{�ື���j5F�Vs�\��c�U�Xв�Sp>T�^��7<.3��L�)��YsI�q^���v�*�]�(p=�K+�6`}�C��(M��fX��1�+�<��2/|¢e'��GN�l���F0��[��iX}ґ���(�T�U��#��_��l/��CN��.��d��#���%c�܇	�<��u��_�8���Pe��)x��mD�;�!	(�5�=Ϊ�Kn�_e�;C0$�솭��Ṯ��q�J:Z��r��B����b��5]9<�OD��}03HL�b�R��5&jo� 5Zh�۶T%}p�F�qW���'=���:1��)d%��-�^SG�\f��G��c����(ʉPكm�H����C�̏�w�&�^�<��a�R�"�]~�� ����w��ݘV��=���_�)_ �4��`�M)qU¶���f����<k��G��0��o)�TM�l@H6��%o|��/}L}]8�BZ�d��̱xCN�ȕ/��,6�3�IH��<���ţC�?m,+]q�x�7h��`�W�O�M���y��)#\	4L�]��2��8�ڱݸ��R�("�c��`yO��e�E����7�z�.V���Q�<߳:P�����%:��dE�mbG����?��L�T��_]��mb h��%+Ww��V��������`R	u�Q���ВSl�]�A� ?�X�8jo�!������{����Tf�J��gX	;(u{є$G��;��?n�㮰�S^;n�\�n��Q�{��r1��q�S0���Șӑ�b���Z��v�ω38�. =G10;϶����_< 
�c4q����c�a�[6?���<�2q�v�zH�󁤪��Ř��u�r��}�F�ƽ)jf�.e��!��Iq�;@ys�@^G���}x;BL.��Q�����(�P�
��\�֏#������^��!�:��.:�@<��k�~��]�F��[�=��f3+����2��I6����^4.�U��4�r]3-��Y.QNsa�9x�jתI���p���H�&qIk�� d�L3Q���W�z\���1�{[J��L���M���šTΌ�uxB�'���o&���h�P�U#cds��u���ʂ@}[�h�곺<j;}�)t&�K/5=y� ۍT��z����4hd*���f�a�SC�<��"o��ɐ=�Z��f�o��Q�+��=)�'�"O����(e���P�'�+���Z��ʂ+��A�EV3� ��,����z��uV����ݜ���u1H#�����Z�F��ky+��@w��Ip9�wlE����r�Ϥ�j�?l����=�:��i �"���!�E�,4�� ������qk�5֩~痶5�$"����w!vo�:ۻ$5Xy�wH��R��#�@y�j�������*Cv6Z~	��k�����-�y
�,��'�DYd�uM,�|*�xcc����Q�W8U�~<�����2�5���pWM���r�!��lTL0:��6":��,(?�_?�)pL�{u���R���KK:d��6gX,����dN���>Fhě'�6!Q�.�r�˜��u��L���=��o�䣭�ש�X���B\�>e4C�k}��N 7��h~�:�M)���ĝ���l�"�,+�Կ��� %����bO^W���s��G��]gK�vo�3e�EE�ӻ��`����䓟ў�OۤLQ�q%y���u���ʕ.֥�Ҳ��R���JT��q����UA.�sf~�(��G�	c��qtL�2�B���2�I��E�B�"��7������m��H=�w��R�);	>
7�/��S�t5i:�]=U�	��r�'���VD�A��J�C,��`�J��2Ѯ��m����r����fiq�)U���b Zr+b�nC��tf��*̓4���0��J8�aŰr����P1G��ċ<�_�3xm�8�j
$!d �q,�L*]q	�B�lʜ���;�+	�� �b4�	F��>�C����w��7N"��7QZ\��#yIN��a'*���)>~�����y1�X��)����MYl�:
-b�v�t��>e��_\���S��|�vF�5���DM���z�K_��l!-���(E���di�;��K������?�5��Q/3[�R�����8������BB��]������f4kSk�m��N�wyqq��f���K�0M�E�3ˉ�Jk��B-(@Zv���W�x�ѿ�9=ɺ�6��( p\�=< C�$���Ɩ��4j ]r9Ӯ�?���5-���r�qs�
���g!nK3����,u���bn��H����"s�8�^���l��
�pr	U�����s�g�ɷ�C�`_�	j�d�ٷ��_^Ս��V�����a���X\�)�-��K�O�Сq��T���-`
Ȟ�����Zq��x���%�} /o��#\���K��U�{�pU>�ۥ�`��#
�o�pmt�J�t��� Ȏg
j{��b�����<ߤZ(�xB����>��6|���[:������Ŋ4��Z`�G{�w�>_�h��K�N����X�J���sxD�����	���yH��#\4V�k&�gW)o�	��<'�4^Bc'��+��<��F�}o��qIߝa�UK Yz+���e���� J��T��+c��/C����� hր���J:k;��=�9�ٻBN�?W�d�B:���,A��%�;�VL
�þJ$�:��2Vp\�o�}�%�j�ו{h�f �?5����4�7��|���db'��
r���~�)z�)^�%J�f|h�6+G���.�kf�{����տ���Xi	rŽi�Vmnd���2�Wܿ���0A,o�p<��Z��6."8���ۼh��-�m�e�*�@�eĲ6y���(7�q@�{_$P)�2)IYi�oPo^���B_�idy�f�_��0��e %�ۆ����l��Ed�q
��1T|ͬt�?ɝ��d�6$Ҏ=�N�3O��HF�X�Uͧ��,!��AF�q.O����0�4N�G��jy���IЖ�슑ʧ���k��������$�C���kz�Xj���$X9$�M����}� <4��P����c��+�T[hj$1M \~��D?��׹��ZW�������7{ @`Q��{}-5l}��;gQ}i��sE��O�S�UCq���:,!
"����	
���#���{��
�&��2q�'k�59qPC��#��鋑D~�:B&�O��l�=W�vg<;�d�|�^I���e{�}jh�+�ˊ���hy$pG[+�Hٰ?գ��I�2�qP���0l5ޅ�В���2�{n����$hڮn�}�j�T�t~�'�>Bk�B:����-�""�����d��VCΆ���a�h�1uo�@$["�Q �+����ǂ����?� �O%�q�Nr�k�	�T���%��RS����O�����$�J�i�B���h��O�m�pS5�!��>��yLU��èTh4��Sk(��iEC��`>�nz�����e��B�-6	��A��)�ӾZ���j��zk{��gn����@!��*�Z<f��(�y'�N}c�*�m]X
�=����׍2uDw�m"Bv�Su��(H��۾]2w��� ����6Dj�����	�N��z�G?;�BX���rJc����`�����P�Y�i��9j�{��9q���Ɔ��e�Y��K�~evt
�N�[�h�w��^X�0x-�l̋���X�.{���:@�Vɍ�$�����z<�6	F�hJ�ºg}D'����<Q ���@�/}mz�ה᎝Wù�4<����ޖ��E���VӧH�C�^�e)�v����j�96 &�*E�ʳ��k��gG���H�c�e�Ь�����4�5��rQ0K0�kj��f!��U�'$��`�%��.�Dr%22ק��U:��h�%�-'�j0P��W��wF�:P�]�P "�}�ک�M?#w�������S�=�!-���Y�d�"�M�c�yL���*A=7il(�^M}�Cj���.>��37��ݱ��դ��B��Mجt�&KMG/8@����'�T@�uM�L/"#4s�:�BkD���t�I(TP�6,:�/����R������J&7ָJ�59h@��ήaI�Cx���4���&o����Sl�>F�D����N2�?���_:���u�{2�\؞/]:6н�3#�e�S��	�g}g�Y.$3UW/�-v�:Y�Dߢu��\ �Kjd`�֡o��Q�u��:���E�[h2��~�^�oP��ӛ��5f�b�ds��h}�@{ts�ƕ����z/��.�����9-�+�	���4i�+wG;�KVG���7mv4�c�E�p]���uA�����d�W��k�D����z�
�4PۜP˫Q7o�A�K�<�����u�ΰߎ`���: �^"��3ٲ�2<T�`V✷*�!����l��G(S��"�����N8���\�BlUY��@^E��k%� ҵIC/Ч��o���1�=�7-t�������X�{��k����^}u��=�A��P^�����p�k �b��{�/�)��Y��6��B�p{���cאo���~�i�:&@�2�7YY��浃�%5���ۼá=�	�� ������f�s�>,�J��5�OK������=���`on��o�7Vk!�ץ�=�_�D�7L#����0�ȝ�ݸ�P"�!��#<���>� ��M0N(V��`/��¡oY;�m�$�m�{��<jt|a�N���=�����eE9J�o����u��Gޥ&l�5Ձ�)!}9ۚ���NDE9[�'US�
"g�
v���4E��X�8�X����Jߎ(V?����_ ��v,1@'J7~&1����9�s�A�$���
�!�r��"�1T]��#ZL�1s/@vyA����wS�z}aʋ=�BA���8�f��''���~��0K�_�E`�'����捃Ԡ�G����+�m#A�Yr��쁷�o;ClG�N�*-kj����6�� �8̋Q� �6��"��G�Ȓ��R�ΑD\�M ����rKM~A��oI���$gE��*AO�į�O&��\�i�Q?sC���;Þ��M�X�^��t[Kл�eN.p7o���i,߼CN:F�H���}?^@0-�@5la-r~���QGg����N������;�?e���!����R ��*�;��첥�C~ӑ�'�K�� Q��z�G���,��Oj��*|w��,Ie�xT�¥ֈ��i(f�֮��������s��!%&��hvD�θ��L�Z�Hi�Q��l�6jVW]Iv������1 ~7�{#؄��9����1�i��M.�k�\�10*���ӿozs&l����&���Ą[F)�f%ť(՝U�>�%�`t�ڄ�~P:CB����e#׈�H��9�a&�Z$CK䬔�-��YF����t�a�Ug��n�_>ʋ���I�Rlc��H�]�	] X��|��RͷV`�b'�\`�Ǎ�~��1����m�9���ʩ>��������c����㒷� �?+��9��z�*V�K�`��k����}��E��ʎzT�"�7��E��sQ� �̞ٝ���(!oCc���`��:7���'�J՛3	�?�f�յo	�\��f�Z+�1����/y��r�����Z>�W]�9����N!z��7�2 ����cWKmo.��%CWb�`_�["�W%;���+��{���u�?��O�&]�zDr<.6�PV��l�0C��.��$�G� ����F�y�5VIQ:�Y��q��	�f�v�>��:�ԯ]��lc��y����L9,�@��ݼgu��l����̳Ӝ7�Wɓ@�Hw�����	�Pg
3���He4blZu�u��͗6|��c���a��nX��=��2��e�q�([7j�8c��$A�{;�.�&:O摋.:���Sfo �}8,;��qm��|�-��н>�՞�H��N�������*��3�Pvi��*���D�1�zQ�w�[.�-�p����l"��d7Pb5�� �\�-2̽�I��d;�g@HF�7ܭ�$��/���a��G[�k�U��@�j�vrp2�3�'VV�oLu�͎���5�F*���+���bC?�!��"
4�%�`b�Z�P��5hrH�u=دE�w��;rd@�����:Jj����]{�k��s�닎Cs�+ɳB���>�J�+�ɰ~N�|?�k�:I꼒SZcz��H,Ys�]���~�m����W��yRd���ٲ�uyp�U�EN��AcA�Y �;��>��2=��`�H��.AO-L�l�ok�=�,0���w��8���e�.��{�}�$��bt�g�''�2K�'�ހ�^k��o��WH��Z܂Ǘ��¶����$��t��B�� �!�ջ��KsVp�u�����(d��r�)3lh������g���]���胓Jus8���޳�pG��#���m���M���3���Cx}��g�;o{�����?ٜ�����Έi 3{5}�DE���6�5h>Y�D���)m~|5+}�Y:�jZV��9䶳8����E�P9h�ٺ�,�H�D�yp�a�������.�7�S4�G��#����۠GK[�1�`��G���̇�3���W��­�Ƈ�6+_������
�<g�AU�(�H�`��c�V�4V�I�IX�~fB/u&	�Ӫ5b�
Z�A�',��
��b�>_�{��ݏG��T�fh�wg�P  �z�R�V�ݤ҅o%��6ۈ�v��z���w���ґ� �9	��v�ɠ�D�����|\�3m��[jC<؇\lO������q��.�3ߔ����u��oy��)�N�|��fP<1W��~oxIl��b�	Pp�J0��B���[b��]%�<����W��5NtAȫ�w���5��p}}ɍ��OEQ�%�p;T�p���wU����j����H�3݆�?S��el+-�Z4�#r�Τ(����2i��A��>��\��~�����C�#9Ly�pi*�uӎ�-��q��¸*-7����?)RY�iO>m�A�6ď���+�3
T������ˬ��N01ʻY�&�gV�_��L48�S"�|HU�;��.�q��-���5�٥��N-ĄU�KB�1Z�Z�b7����Z�r�L?���.ӓ�`�&g�Hr�&���>�G���
Yo�d8[�
�Y���cTQ��w��策��;���P�����J�C��!}X Z�Xt\��,
�b�G�*J,�^�&pd�]Lm?MP}����3�/RϿ��*Gʥ>�9 �\ְ��e{[�P��p���G�p#�T�a�(C�^A�x8��v�L{�)�GF�3!G���=���)X����l�퇂��W/ˉN��$���O��C2���Ba��������F�ih�x��?��(�|�l�dD�a���;`q�>QR
A�R��fP3�J��6�|L<�J9/"~�r
���/J��!���U�I:V�H qŷ����뼙�S)6^�GO]S�������t&=*3X*A�cwz�DQm��"h.�i���/�_�r�<iFn�(T�H	�6�5
 D]h|=�SLlsQ���ʈ��`΁E�ʍ���"'�8�Z�Z_�w��e��4��OP����ua4��:e1�d���T�e�e���^,E|eQ#���Z�d�Jg,5w�)�ڤ�-�Na>ִ����%�ւ� ܐ��M&� z^��n^�]/�usԻZZ��ūo�v�*�#4/�A"\`�M��������*Nn^�F2�t�4P��~D��QoB�m���.m)+�Q��2Cu��썭 �b:X��?��0%���ynL�:;ӟ|�=į��]ᏬeK��l@:I2�J4=��a�����d;��p�~��>��v��^�eqp�����gv�����mh�ݢ�����wӒ�Y�M ��#�҇f^z����U�{F�p=*��eIzX��D�*��[׷
	�J3�>�@�	�2�.�M�&�Rx�ۙs�[���t?T�De�d����	���ʀz^�_U��v����x��Q�Z8�4&�)����MG�hc������V_��������8��.O��Ӣ���)��w�pEi?B��,�[�+n���4�\�d\�s�1���k��W��
�<���aA&a��e�ޢ�2���h��l��j����l.!�U[s�s�GV�ڶ����v=�X#77VR�1Th鐈$7���=*�Q�H�$O��M�ĺ* �BX]�C|_�a��x�pGЀ�{h����7����+d�~��
�)��^Aյ�@��4,�wQ�/��SSъ]��I�-]h�K�������Y�^��J�K֨��7)�bl~񢸥dzB�Oﷅ� ,v��(j��7T���=+�\�����$�%��I�q�]|����k�06��	����0����\4c����%*�md�C����'N_Zy��]��}$*يu���Lv���X]�l�(�0D� �����i��� 9�q�.6i+��<f>�����?.��l��Dh<�DW]gd�[�Q�t]X`��Ԧ��ʿ�U�o�<ĉ����)�m�̃7v�	p%�<>�,����C#K)��Z���Jb�S2Dw2���@�(&�`�#9���h�P<��@U;�k*h�d��p������҈ʯDӦ䕤RE!���}FE�Os�x�I�	UE2Q�M15�(6�#������;l�[������c�S��/8 ��U�n�cm�W���f��9ww1k��� �i�rl���t�����ntw��f�x���"�BY�9Ǚr���;�0F��&� 2�0^ҥ��-��]}' ����r�3hLQ�y�.b�z�V$*�,W"'ӭy��AGh`�y�����," ?�_R�A�4_�G���6|�� �y�����:��_�(;�T�I�P��^3�u��.G������t���m�zCOve����['�[i�c���x&�íݷ�<3� "H���"v�c��]��e���W:W`�;kW����8�F�8U���=�-b�,�r�T��)�dIx�8�un"��7�1��+��]�m� f'��W�;�-aQt���OvNM��z�f����q�7v�ߘ�w�ax@�ݎ�Z�e����oiB�L1�7q��V�5�Xx(�ɵ��}�r����-��.�� �K�����n�s����M�)>�s�~x!����S�ѭ��̆S�����Tz�쟠������ky,;ŠDq��b�E;�_B���E�z��1��;�[���P�؆�Z}O�㡖����[VR���ة$�N����֘� Z*�hӨM�ïJ a������B��<A]W�r����UP��"��b��Y4�{K�il�j���Rڠ�*Axd{pv�o�;��+���[��c��J���G-�k�`&K��|@����x��evҥ�&��r�"60PLj��/�U+�	�h�i��:��:~���?ce!䁃k�1������n
_TV:�.�
_�*� ��V���YO|A���;��͆��C��{�[B�ݴ~z8���.Ÿ���k�9\�pOu����W��UEn��6��/��\��������\h�Q��x�gi3Ĩd����V���� �|��?dEs�HlC�q��	�6�8�@�dAl��P�
L2��W��5���Z��ĝ	�k�~SK��m�ԫ��{����ć˟Y�o�ԇ"���� �ݪ-n�X7�ߟ���5���Av3?��8p�V��AT��8iz��K����Y�� ��P�O�f�uL�K��Z
Gd�"b����<�%�����0�����	��"QRX�1��D��QԤ�>7��쩋 �D':j�G�sz��+���@��-*�K�������:�ù!1S�+2Z�Jp=Z���l (��>�űG\Ɔ����[ᡱ�2ni�'|�'7t�ڠ��{�u�J.G�XM��Q�!�*���r?]���QH{p��Rpr׀P�y$��	��07��1i�.�$%J��j+�8����Z���Y�f��{r����K���*��χ���3j-��[o(U}�;�y���,zõ	9�J�����aX����ɂ�C_{g����9]����ȟ  ��ϟ���_��y'_�57@���ɝBnY��s��3`��m])��3���ʀ�j|a:�ۍ8DaN�Xm�o"�Y�]D�G�A��g�dc]j��d�!����l]ڗ�g��S��%��f_ԤMˏd�A/���X+LBs��m6�K�?A"ݴs���I ��+?k��n?�� _q�\D�����Q<�'!��\�/����<�i�P#ܭ�HJ0"�f��_fa�ΌwB=�u��D�"w�p= �(�I���&�����*2������@f�5*UA�?�)f�M@1�v:/S�H73����KL��		vH��z!��!{�(�|��U��f���E�-�J%���M�w�p��*q��V�4a�''�S8�PN����q&�]ڼ>u��5��
����/�����_a��!lV3��Sx.�o��[�0�98�k�T[5�x�o�ˇ\!+(쵙�����y�����d�}d>��@�$����xqz�5y�������PS�G���U�Vx)�=�Hkޗ\�uV%�w��ࢥn�7��"1fR�g�j�\��b�P���h���_��;d�(b{�!r-�6�ݰU����tIw�l7�Ҁ�|�@6�<y������9O>��)-��!.^��\��f�!�] �w%u�f^�*�n�oT�7 �f��� bk>��
�mz�f)��"���&�w�2`�2�(�<��;^��� 
�zd�Ha��y�jʃ<���=�XoG��l�������N�Hbm�O���O�Q�?����h���Kh��)Ɠ��h�]����[�/�v�p�h�h ��J(�71�� T�Q\��>X��S�gn@�o������3�x��5%�,��ɓuc��Ŵz���.
S�ᘯr�K������������u���Y"���m^��(�_%�R���9<4��048���zȖFd�&vv�N3�ജ�uV�n~������F����|Ӭ��O�D��)��gy�+�\F����k���/�.�aZ��w�N�!B7��M�YX1\7&���O%-M�ԣ��j����6��G�¯w6��b/����w9��3h27]�kr7����(Xs'�G�@�/�#x�z09u	��;�>�S�<�ܽr2���d��.d��s[_ ���>����͌��b�K��C�y�d���<��>\�T��*<#5�U~F�rB�t��C-}�Ezb,�dݹ�����f�3P�����ve�YM�)l��"���V�i-�l�������j�� ��(1'��F�']ӻ�$~t�e3��8�L�����.��YHF���J�����z�BD�Xq�hڤ)?�M����G�^�ݢ9�QxXtPL�Y�H)���&��B ©�X��%|.�R/6�`D{#׻L�ֻ�F��(���#"�b������U��:���Q���?�ًVLV6,���;�� ���G^���99�QӉ.�a�~罕9E;��`N���C�{&��z��
�5��$�7Χl���M���M�>rm�o՘����l(��0Q�\70��H&��O�Nu�lL�h�5�L���������]\Х�yFCӕ��}n�vș�|f�KG������6,�<։���~�c����yC��I���-<�4 P��� $̺)�Vʙ5U(:�8P}�����hL�����p��xN[�<�7vAh���H��u��3`sC������B(R[���Fy�GE��lW�kQ4�5��q;Ho��f�囦�|��P�AD�k#;����B��銰��}�$MOZ��$uhz����&�� ��s��� L(��R�p&'U�k������c����2��Ĺ��d���ğ��9�ez{��ғF �,���(Y�՟!෤���|�c��(���d�#:��\�:�{���ג�7��S'�9�`f\)�O��KL�M���i�ܾ���CX������!zް�؄1�b¯�?��K�}Bi|�X��XP��y�t�T�x�n�Ϧ���
 9XA-�a|.���g�OY6Mp3��Tp"��f�VC�O�b萧g2�GY'��\�~���TEa�O݉����Һ�k��8zzr!�e��L$�[0�������*��Z���)����>�cGٓ���P�ZE~��>J���E� K�5�8*�'�H)�jT�Zf�k�J�����U*�lg'L��[�Lhk�r�IH:��pdKD����8�o�8^��������[QE��h�hDL��Fv�D�ű�P�O
� A��Dɀ\S��"�MX����0��1�PàЉ�'B����N�{��a�W����Q�)F�)A;IZU�dc��q��?"�[����q�d�h���V
�d�<n]��5�7i\���.Č;���;�#f)��q;s��\sE�r���#��2E&(0!J%7��N�Ի=����kl�c�I'�Y���~Hdwg��� 9���f��o-��)����co����Z��藍�L}�	(}�D��:�����75��12�l��$��a)ʔ?Բk*�Ž+>J�7k�r2�cNNT�U)��\���c>.�)J��
ł�nI�aB*]�(H'y'�F���X����w^���e_��v��Fg�R��S���{��q��˨�Xj��P�J$��0C3u��� �ؾ2���2�6�����j���K�RD~�[���3+�9B*�)�M�x�#^%+�����#c/��ݖ|'9+~n�.a3��FONp����%��)�码���j,�	�SzZ���-���l���#ǭ�h9�K\A�୒��|������Tq8]W�����0�5�G���|dW���G{�+d�i� .�l0�ݣ��H��Dߢ;O��?k��b� ��
���Gu�*f�tn��귥�{�l�33�_�A�}����ɏ�x
#vb'Hn3�s�*ڷ:��*�Nk����8O��ҧ���H��� �Ȳ��,��?�Ax�O�Ï�%d��	8�|����ݤ��tX�6�MTZ.:9vW/�^�&�Ň���]�����ܴ*��r<����ķ-k��� o�8���
���eB�G%�S��/>�3`�-���;��<�(k�lC�08�i(e�r{���NJsl��(XkQ�f����E��/ʚ��iX0���Ngu�IҪd�JY���d�������鴩	�r��
�^���� ���Ƿx���@�rζ�)K���@���æ,���t���.�7�݃d~n%�[>�V��J�HG�\q?��=������S%��ǯ����N�C}M���r浅dx�m{��
��D��6L�>��D���܉֍������VoN�v��C�� i,�яC��a�Ѳ�<�; ʏ�i����tt���b���{��8"���������� ��~둡�135̀�poN$Lkֽ�c��o�7����KJ�^rJ�K���,l<��d%t��8?*�JRty�~PtT���V�À��H%�n�Y����!�0[�>3S�Um����hb�$p���;[T�	YF5�����8YW�:�����=���1H�Ubݍ��lw������jɤ�q%�su�T�}�Ot��IϘ����8;&�M����"-�����=�c��L�,p	z�`�8k��8x8� �N�R�m�Y����>�ó�}��)����K��Mj����Ox;ݿ���Hד�����e��������#�6�(�J����K�t���>��_.3�T5����4�^r��ӬD!Pd�����Z5�Yv���5�Zc� ������JǼ@G�������>F��K5->����s`�D�;���`����Pǹ%N���~':�
!���E�=c�FD^9�g���Ss����%����G�r�{Đ3K3~u�ܷ�ۨJe�� W?`������E�s�ZW��'��I�j�Q�VU��
T�?�P�>&�+��g�Ƶ��#'�9gio&[��*��J����O�dS�����b��8��w�sgi}x]���0��x�V�B��aK��qZ�T�ux������ʇa��|���,xڙWZ&:��f��SAu}�x�R�~�|��nt��Z3u��xs��0��&?��u؟ՖԿ9Ѧ��M��Q$&��6R6Q�o:GE����k���������FT�9��2��Ӆ[�(�2�ą�a4�R9H�T��Xe)/���4>���{�ҫ�7�a�����X��\�����A�,ԕ�T�����]��VZXT��̙�kB;9	���[a3����*+D��+�������:��C(�\,�
��p�e��2��3��	�F%9�@F��*n���WB#
xx@��*��� /X�+�L���`7f+o_��3�=	`�*�YҐq���{�<��/��m0�|b2��	&��?�[a�I|ϭU�Vt�ZF���漨�x���L�Iw<Ȗ�C_QY��<��p��&�����&� ^O�93�gԗdvK�=�J�N�,����#!'���MJ&��~8��$No+��1�����KBOگ�j�x�1�V��h� 'f|_�W��̬���jk�=AT��[k��+����ĎĆ��Xe��$������5��a���TT�N���L;r	�?���&�~`����@�	�6"9"Ys[���*QO[��f�"
��"�"�9�`�����}��#F�����}�2A:|-Æ/	����$5�#�!5ě���T3�yd�;��9>g��؀]>��g/�%İ��\땙��]��e�C`����m� d�h���6,v��!ݙ~�[�L��}$�y+_���^k���Zf�׵�_��D���GҬ�]�S쟴-	s4�٠��������$qҍ-fEI�d�H�^��J����:�)���V�ի0��p�2��j�a��e�=�e����B@��an�����it�}�'׳���5J+:�(��Z��^Ԁ�㤝��m��Y��>�s��,���{����:Є b8��A�$'��{w�fB#�v����zE��Z���_7?	���vN��g���a���Y�>^�������",�޳9�l�{O��ߊ��cT2�l��:*��#(�T ���4`��،��K*���|0�I^��l�%���&����u�B2��F'@@|���fw?��~�=�zZ!J�J6
붃�r0��W����/�%΢G���ɒ�J�V�gk涅wN�Q������U��|�,���	��S��dZt��4�9����{4%�O����X�z���9Z�N�	1y�Ì��
`J{5������I�p#LU�k��S��k⌒%Izؕ�X����>@�t�zR�E6���:5�k�
`h=���������B�l^���=a�EO�ڭ�Hǥ��~[&0g�nѮ!V��=�倞D["���Nü�s�*�����, +rh,��Ϻ�5�}�]��l`ɍ�PWo�	�]�����Cb�~�20�X���i���V��>I��4��K���s6ʿ���Rqc]�X�PQ�ˠ����O�%�N�cd���ɔW�a��R����(I�u�-�^nL���Y˶l9�1�t[�Y,36��34�&²�T*8`�zO��t,s��i���c�j\� ¬C\:d�����/����d���������
��	x&��u�ɀ�в��эG�	��uL}�yiv�Ѽ=�_6�3l��s�XGe��"�u�} ��w�hcڱ+��>H�`�ƺ}�"��]�= & ;LlӰ���"V?��Y�dᏼ���Z�@����7���B��Lx�=.6�týyo��ӆ�{<V��Ђʛ�wb�גjsS?���ȗ��>���[���e�XFИ��"����e[�[o�"-^�H=���*�R��jkWɩ���e"���v�A���Z���φC]`3����4^%��X{�.A�:Ҕc��K>W�K���!�ZJ��Z�is���`��d,Z3�Q0�|N4�����V˕N3��x�b��l2� .ӧ�u�����D��=�?��L���#D���'Dϭy45%y��n�4���,C��$�����6��xB>dr��K9�NGG/��u�N�r�O��?�Xz]�0E�m�G��۶=���iÎ+��{��a��1R(K�&����!���h]�I�y�RFZ?��l�;��A�����|R�v9DE���={�b���Z�xD�(���^j���!~y�Z)��R���H\צ��݉D./�:�Iں�o��5��,�o,��C��=d���S
C�D2G4h|C3�>v��|k6�.�>пC(F^8�1tF�?��z�c��D�J�?��Vt�L�_<b���=6U\�RȢ�	+X]��fQ;���J$o��Ѡ���e�&� �巳�A��n;��ᤣ!`��3��׾����}C�X���������r�E|H�5��\��Z�r��U�`N���㟐���C�c�-eog�~�������E� �GX �i)ݩY�?�%�K:���t��G
�Iat�Ȳ�2;ԑ�ڣ�]>
�9�+<���<w���-%��Ƒ����GZ�U;�YT�B��%*����d��9K26ï��]�A��f8=�t�Q�iG,?<\J��(iwjq[�k�l+�X���_�GK}.$��:d�zQ.߬�֜�����I�ח�q� ��!�]�n����t�h����*J�k�k���j�hŀޣS"���.:�}0��3��2~;[ ���2T>�`.{ň|�� &�_�?a^ʁ�����A:��Wd��%|OR�}�3Г�&�N�F��j �Qpr7��/�?0/o�e����C����A�{f����Vnd��Ô�.������umݑ�ϟW�Y���]�H�*�Ñ~�.�������,\,V�!��(����Ő�y;�P��$5	-�����$�d��)�����j}��IӜ���s	���U�������f��KdS�Z��g�'U7���$�ƒ��sqj����+�m�ļ�LfdF��*΄��24�׋8��+oP�޳��/��(>�?w�LRR;<���]`u ��S(sy�i����8�=��D4���l�*���tw���輡G˾���.��v�cYp��k�j���%W����\O[,l1y�������**��_џ).�����2�O����� tY�9KV9�)��l0�kE�����M���������[�@yW���y�@Y[ì��h�<8�6�L��5��>��c�9\%�F�4>:Xl�5AD��������x�2�'M��c)kSk��~�Ou3����6���{�1�{���7�g8r#F!^�Hm�4ѓ�lG3�WO!�
4b�G9|�1�΅V�l8��[	Y��ʺ��ޢ���!P=�F�k=4�5�$��Gn3j�˧ي����(mkԳwۏ?W@Bj�In����m��^D������k�2�Ԗx~f��	�G��m��,˶��s�'�<Cu�T"��ؚ9��/�H�۷rXW��lޣ�Cg RqJ��$ ��v�a6*�r�t�q9a'tW�ۗ�TX�4H&C��i��P!��0M��2��e1��#�-QP�,Ik����:�R� *�.(p�Ø�q��qs�Rÿ�����'oS�4��8�i�P!B&R��x���($-*�L��k}�8؍s5��a��W`��T$�Z���)���mb����t�Z�����-��� �Z�%�_���7X�(���0���n�. �V�7RԱ��a��M�� _h��/J�L C��~���^��b9�^�'�������9�Qr����)���0�V�(ntL �z,s�7�����\�� ����t�f���Ͳ(~�fm�j��d��jA�SJ�����E[8ƀUv��Mc���5s+�utI�6��
�X�غ�/&a;l��1mb�����^UGz-�Q��F�BXUf�'��H�}J2f�y؟`���6��D|��+�U>Գ���[jh��LN��8�5&=3��v}�m�IYԦ�-!��� �v���HQW�:�,�P���!��v�Y�c#����d�h؏5!O�>6	���w
��h��A���]7��[h����e��V��e���4H�	O;���c�r>�F��j��(�wc��p��Q��hSy�ٿ�b4�ڙ�	�C�Dΰ�>,1�(v� �aw%]�iU�k3���gzˠnRכ��<.�Ó2�VS��β�m��쮙D�:qS��B��H���ɍ~+�|���W|�ц!�Ȕş�>��
�҇���=+,�3������s �)B�r����}��5A�d=���TB�Y6�z+�N޸zESr����-}�`kK��M����b>������PU��K7����E�u�툅"�J3� �R)���4��(^+g=��i��W�X�H]MǯߎΧ�{IX�qפ�H���Y7�+K��ܕDmE*�|�w������o�q-,|we�Fv�z��` l��'Ɍ�G��V��Ik7��2�@�̓�,����UV@�ɢ��Q����J�lgb�[� p�%�	�E�H���Q�׍�;U�v�S�
��m��K=4�,�b	)�Ğ��,MU-m��n�K����q�֜�;������h��|HS���>f�A����4�6���;R���U��K!��D�}ϰf�F��7Z&��!;h�h����n��j�}R�-�m���4��S�^�"�y:߲������
�j�J>k�&Y}���A�O	PX-l�/�RB�����۬�5=VPT��lo3��F�"n��P�|Fx�i���:���dݢ����[��ss�=xj�;Gcȫ4F4�Ї
�E9b|9���΋��nFH8�	�/��-m	�{������dP��T�q�v���������yê�A�v�x�&?�I�#���p�#|!����Y��2��
�rm�"�E���֑�p���ws���#9l���z�����
��*?�Jo�Sn�D͇~deO�������1T/�N��͋b�=��i��Ya�sE��2�X'�ő�&���-�3�_�k2���Z$e�@}��Y�R����(�-�l�(B59�Xq ��@��9�n_�{� ��e��$�b��闢����\�޻"��RߪB�k�5X�`<����3������X}�s4K���u�r�Pg��fwIT��P�N (gb!�pl��rMש�����w��R�v[�� Qn;\"�`���7��Ȋ�Pr���ɀ�	�t�S���BȤ-$��c]�k�6W�a�mC�V�}�V����{x��m���P��\W&�(��J7
�iSI,��*+�!=��:�U-��3��,���ؖd�U�N�c�3T��
��#n&��E�j%ܔ��u�l���4�s:H,��G0���~'�[����o>9I���(����S����lv�H�:|���r=`pu�se{� =.�r����aGT�̦Ρt:�����G_.Dh�:����W\��:?[�U֋��`���5�Z��-�G&��a���'2헨*Et	����&���J�9���n���h;t?�bJ�( �*�L4��6��+�ͭ~Kӣ*_�К��՗enjG�ݰ��'+�?9
��	���uJ�yY/�Qj�U�v�*|�h�������o"�>=������d�� �P" ����u�Ì����nE�z0�?�2B�O�'��C�f�+9Q*7v���'P:�TK�m����1�g�;��Q]\9�,��M��+��T��A������d��՗u��o=p�S1`����c�F_�Լ��J����M�=(,���/!������)I-�+�mk_}�r��	���I�FN�_�[�2�l#�Ě%���`<?���M�_�$��8ũ�[uZq�q��.�	S=�u�j��\-�H�,w��6)oj�H���� e��w&t쬳�(��0��eL�_^!��y��-P#�3 ���FN�a5 ��#6tjV�a.���cVPt��dT�}6<�`�P�������{��9z4U7g��1 �m�r���W.]�]�j9�c���jٽ����R������S*�Ab����Wz��c�	�d��
�wb�&�f�ꝏc��O���`�ߢ��r����^PhDIq�\���T�2�@�(N�r.�����VC�	[��<$�#WH�2@� �E䗉cJ�9�����rF£�EЉw��}���C��3%X�V�o�9|S�.�s�%����Y�ek-�g���K�OR�{�������XAk5�1��QP6�12�_a�.�E��H;$���7"���YQ�O�ŅuR���� ������Ka�����7�2\ހM�`���b-u�6$�n������i�1�B�Cv#��o��#����4��'}��9H �9�0V�gM���Ҕ�d"tغ�0)n�Mv����"�Rt,�H����+��d�Ӗg��կ��}����B¼�Wa�Y�� {*쨧L�Oϊ�𞮌��Q�I{
� ����3:��������k%9A(pdz֙�16ANo�����ADYc0��ow�K�&F�*� Gok.�V5x�du����[|Uk~���	o%��p��zNꐑ{��EP�i%�I�Vm���x��0��Q�r�Q�O_����pU�q�R�*`�2a墍��kb�i\��������l�����{&������ꠦnW�w:�-���6o�ni�-��&����!Q����荨�²��o��o!_Q�˭�)����	y?��OG�K�s�����<&����x��d#����2GǢB-@�LeOl}���n����A"<Ͼ@T�B<�:�{1��g�O�q6	�7��0�6�m�U�FYd<7�=mڶ�yMh_�9�g5T&�'���,��\Ư޲�6��pC�)�Z���jlv��ڵ$'��� �F�#�JR���J�ݨk�\*H��>�2�-����=1�ok|y[ҶN�z6by�ػ�Y%���]u�3�����6,���w���	BP9��Jj��L��=�y�8�;A�f��;�[a"F)�]��VT4$�g��b�X.i٣i{X�[:�^���[�#��Q��**����|$�E
��,�\��@��
�\>�=��8������C\�u
�c���~����#3O��s�={UGwۇt�#~�6Ud&�6j�Je���l�0�+�<�,+J/���0���PE�!5	2g M1�E�5����(Ꝥz�n��4w��0y��M$�,R�����fuy�D��6ъ�\�M� �Z��|5�w:0bkLY�:]�H4b�]O,'�dU+QB%�W�fJ��:+�Q%��:�Oz��i�3��t<����Z���KD��RJ�r�g�8;ؚ����b5�$<=��X�"��=\N���QW���bg��ŝ�2��#|S�S=�ǃֶ��|¿���
���>7¹�u5jlVj�Ϋ+�m�T���Jթ�Ɗ��N߁�8�l��eJe�������Bӛ�[�ր�>�tmű��f>P�Um�e�}+���[:������.`H�p^�>�?�C��Lt�䰪�|@���N^8��
̢n�~N7�g�E���O�^NL�agR�$��\�r\Fy�Z���f����k���aô���Ay��tY�E�79�����ɼ�#��t�)m�	�ݵ�i�u�m?��߼R��������Ja��&�cY�y`,�?��V�8���.j��Go�s�*���6���8�@hjY6��g��6)���b'�#��}Cp��
/��2�μ8�95�4�,.N�K#���	/Y�?+��*�LH�_9d>�I+0��5qgT~�V�|gL�LoP@���a��Wg���Y�s��瘽ѻ��*�fRW�W�ï[,KH��(�ПS����8���"�+���`ɦ�z�e�$M�ߖ����ZB��W����0�6��6I��T�7���*6�5y�����U��Y�7rj�9��4P����p��H%����i��U�ϯәAJ�C�Fm�&����sa���e�`�������)R\﷦��'&z��w��WI�L��+�3��ͬ)���dG���u������	��]oO�Ѱ�0�b	&�mց5!N�J6W57��I_�1��̩:�1N���O��΅L��H���c��iU�?�F�99�K�w�#�#���NI=`cؚ]�#�:��R��4."�� � x�?J�JV*��!&^I-�79%*�=⋟�����s�<꼓&���5hw�E�Y�"sQ�+��0K���H���n�?�\8���N��#`#W�|��<"1ƙj؉eI�2�{��6�rBRL�)�>�а��2�D��C<&� 
�;�����4@�g��M��dI��gs���L� ��MS�Ӹ^?(���^��6�/V�Vf3�����ru^�(�P��	iD��Z�MJ�v�V5��ڸ8����	��տ1:#�-e,�\��Kkf��(����"^@��a/7��6�7�r;�Ծ��[[�}�9WՅ��Xl�,"��q9���J?�mGD>�����/�'9o*%����KnY��m�2��o�UK��諻���|+5��
���� ����;\_oC{�Fha\L������*�eH����g�{̸�bo�i �CYj+�P�*W-v�bc>��uR�OLv��N�U�R�"��i	��A�f�IȖ�gCI�0q���4��܈�Dֻ��������C&i8F��%R$��CfK���gd9�ћ�Y`a�{���ӂt]x�f�oy5�Ҹe����,M/:F�Q�V��c�CWN�o>�S�\N���n����㌂dg
�} Q��!vxJ�}i�p�?��ɏ���?�,`�^Ă����o0�5�!l��u~��n��,�/NN��g�L7�ȋ�4)t�sa:�A֩��ԓD=�v�w�P�O�K�|c�Rʑٻ/����������}٪T��\,�Y=�B�A?,�F0a몘fNs�OcɆf�[�~��W� vU��#�9���Qh�c��L5��!�Tn'k1��R7|�~X%bz{'�d4����yp����@��Bj�ś��k��RB�np�l4���iϥ��$[_����w1=F��X=o��:���ػA7�*��wf��T�ұR��}]�2��r�b38��Am�/+D��f���[dP\?\�˱��=��4/L^F9^_*�<;�H���.��c����5��<sc*gP���e����b�/�q��yY���\��� 6�O�^?��'I�2oh"��뤎Z�λ�������A��4\�Z�zYeU��A9���������X'��K�z�y�����,i�-�5Ҹ\zWŷЙ�Q��T���a�+G.mj�
ӐU6�)����wg ��+���~czL`�r���q�#��2��9t���C���$��[0YXh�,J�뚱S��̮Wݩ����J��{���>(:Q �q|,�؜=|y<�������e�e�e��>W����8s|0~���s��3�=����#����v<i#>�o�v�-�
N=��@q�X q��(��}U�9� �|�6���k��Z
v"V�!�(�:4�g�6�O��{�G�����n��˻�6�X3�Fk
b<�^��/tqc���D_e����AW ܁k�0F!��$���k�#��ˍ����P��g���B�����Բj�B H���!�ϱ'iSV����WH=�y4����ⰵu��u|ȳ'�9�p" &�����ol�&�E�>��$��(}�yIݎt��L�;�U��у2�=D_�]e��`.�vo��+�
9�M8�Ȝ!�,_�^�<�k�@x#H�9����Pv���.a�k���Hvi�l�y�@�����Z���gUqY}�a37�zL~xaX�����	r�U�Y6���[o4����zs�)x��v7p��.�&R'5�K�#��X�H^m��*rѮ�(a0Vw�@ADm�<�W��F�@W�w�"�lWQ1܌������G`:��ˌQӗw))�y�����B�1#�/�:*�@JQ����M� l�hu�<1����B֫r���>�8-}��ɏ�@i�o�ea�׌/t���d�W�7�n�(�#�W��\R\��6�����P�E3p��_��B���Vy#3�<Ľ�#�?����G_S+���3��Z?]{��y�8��G,��"� ��y����w�	��6�2S��$؈���g�a`n����0{���c�1���O���p�
��f�x�?s�]����O���4Qn5��6;U�J�e}i����fp_{�/j<Mf�����N�}@�۳�{�T�X�u��'%�����zB����C�1���L�WY�xMC���.�}�`��h�3eEt��S��ި&�T_^6+S��9�/�J�֙�K�&�����U<�F!��-i�#熒vݮ��Ue!�RLN���?aoW/Zk=����K�n�B��ڿ1)㚞az}"����0����Ku��+�*�e��u.�`�9LD�I��a;A�����@�I�5���~v��zl3�4��`\�u!��u�g�s0jD����>1_���,���˿3�� �i�$P��5g�����������π(�T%Q��T�� ��%C��IV��G��w�O���>󩋘���K ���n�{8�%|����=h�㩖g��	"P�`�B��yD�����u�1��D|>�K^�ƿw�o�e&���4��{��6��>0�]�EVc;��4��\�C!uji���[e@�T�$���=����Af5�Y�Ŵ;�V���<�:���r�J.�?�0��b>C�l`�;�ϋ�2aA6!�N��=K��8:��$)��$�:����= �Vp��~���GN���v�q�f�1�w��=���+�EF��$Ip�z��ѭbo"�P'4eĞR�t2��S�+�p<j�H���r2��
���M��V�ćHv�g�p2�� ���c@�&Û�+�w�~�bﯳ��׾���7���Q7r�7�
�B����G��v���H��e���Ր�m��G$�/COX�p���i{��(���������&� �B�������S��=Ǘ�������%exoDm}t�'����_����moT�D����T�aҷ��z�}i�)�L>ºr+�H�
���d�ⷁh&��mlHON� �b��=;���c��hٳ�z���ĕiԄ�UWu}�����m���@@�W�߲k�{��r�*j�]��ҍ��� �*ձ��r��f��|m�/�9�x��>qYv6ws�X7?Ҩ,0��W�����}1[Sa��'ݵ�+�6?��҃�M�x��-I��5�j��h���17���q}aY�S��wD���YZ�q[^���<��*��4r���;���;Ӧ*E8�,�8��r��Eh���A.]�bX��Ѹ�Sd��}�H{��/-p�O )���Vq6��(E$�e�cmg�8}%��V��-�%8�����6���5ր��*w���#�)���Jc�O�H2�"ð�]�{\5����ޫHץ�!��N���Sя����D Q���7"ECn�p��o��ze+�.�o2��4� 9v�5���g6��r3M��