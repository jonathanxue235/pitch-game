��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C��(b�g L�N�W/u��fu�Ȥp��[W��B/�}��`���n<@�>&��jA@N�z|og��(ocZ�[�/'
x�X�$M8��X�9���jlU"Zs���4̪o˿g��i�	`�����*��W*��)�ؾ�����NE�:)����8=�ya~}��'��+a���]L�RH���a�-�f�7�pw�Ts��,�e�����_wĢ�oӬH<�s�oj3}d  ,�J��cfZ�k1�q��U��2���5\\��m��T(�~x���_j�c+�+��5��yb�D"����$4���,�hM�Q���$�ŝYa���s�O.M^"~\�v�Soc�o=rT�F��}��b����ҡ��G@�/�^�(���y[0�xZ�q��7��H=�q�rZ���J������9�4��y,v���ݬY�fu����z�U�=���cfvB�VRh>�X�]/ �rm����K�Ngg�m����3�Ť��y�󨳺���)[�@ܪ���[<��g��U���
�,+����r��w�ALK5�L9T҇(��!�!Zψ�������� �|����O��`���9Ӎ�~ek^�n(��/ě`OX���q�۵���ם?&�pǠ%m���t��|aܞ��7X��P��:4�� f�l=�V�0�@~���L����sR�D�:萣x�]��I�W��_ }����דa�]�M�O4hX����<5`I��\FI����WG�z��m&�XRV��?Ű��:�D"{�Nw�2�P��.�PI~��Z^7�\��W��+�Ҁ��N�id��P�6� ����]��gE��o)�����{��W�����j.�"�./��m���Sͯ�U' ay|�ذR�3J	;e;4?����mL�<�|�'H�Eí��,ɴ^W�L�0|>�MU����C�m��=P�ޒ�zo�Z"m�]a��#s!���rR�\
�;^Tr>��Y=<1w�a���R����0��C�3����VY�ew�{�����H�aR�7A%�]aˮ�'崶����d���T��k,l�$�*��|�4<-�䖨8���I:+DE&V^�҂�d���'�m���"G
��0�zA��E�e�#���rJQ�j�pPm��O����&$����H���5� ��^�$�2�c�#�����e�ֱm��ė��p$��م�T��9j���)E�fJg�)�b��G~)���:V��%Jf~{xzS��?-9��UG �
��.�q��h�������{".>Z9��;r���$������zm�|:�.3�／��	���5�@��0N�I���tc���g�$I؟'�g{'�o�����G�����K*��go]S�����w�"�iq�����yr�����E��W��zQ�"�����V������`�b�I<ǔ)�ޮE_�&u�{b�I�q.�6�+�8�����LUd��Ʃ��Vo����?�����Q�WB�֑�ù�i!p�X����Ѿ�|B �B�i�C�?j��W"����}�0`�^�=�}��Fk�(̜����X��*Qޯ�%�;�{[���엳�}Z����bg�ĭ�t�-T�R�4�M�0�!%Z[QԒ=��v
=B�<Σn��}�s4��P��El���?��W����Beg������É =���Y@��H4�k�0=q4�ba$X����]�z$�P
�?�ϽU]z�pO�G�]�޶ٵr{o?a(�������}�y�#��p}È���6��S�%��3�S��2lQ戵�9o��k�F��}��=��"���E�Y���?q=����UC���k�Y5�mԕ:s��|�� ����7ۛ��H~ũ(�v���Jd�Z�U<3-v���Z���n��9����VS������x��0/�d�*�.���>�3�o���4�t�V�)����Ͱ�q�zv����)#�y�����4WizG\y����S�{XѤo�#C�/y���;�YAӇ�;��N�%�/��$Nyv��u��>��> ��A����6���>CΧA4 *` x��%�2Њ�=(0��~N(�e�E��ێ=�j
�������#aşU��ok��ÄW%�3hG��B�F&�ol�����pu�FD�=;ouZ���	�	f&�l<�٩��&���,'w��_�j�s<%���F*���%gA��u}9n1�0����'K��H��~#�ſ�ޜ�L� �?q�d+�w�Ww��1��څ���X�p���3D�D)�Pس8�:q��S���qvp��ǉ�Hｲ��D��6db�!��Z"g�|ʣ�"KׯtI`����>6���!��v
W��uYY�w�k����gտk��tyf$�
� �)2n%�2���ϲ�B����&R �'�9���t\2d�*'����5<91� qa���A�[����QRl���FAƸ��	5
 ���g��f���Ñ���P��g���*}���E����:V��X��u�r��@���w�o@Sf��n�B�A��P��BL���֘�K�jtBA[!���W��`�FYJ����+y�$�%�������~b"nuY-cQ���O�-r)=�Q��K�~o�"��[�n~�n?��,)����-�n[����g.�P%�ﶓ��f�������4�M��@F8L�[|�#��b{?Y� v}�#�ˆ�/R�e��Œ���]�[G?���@����i?�~w��%M&-�>�Ȗ�@6p�,�Y���ڠ-k�ޒ����A4G����I)}�Ҷg�]�7W`	'��_<��e��9��3�.����M
�t	#oP��V7�iށTL��=�Q)k����!Dd���_YOK�cy��[��Y�&���0�G�	��c�o�s���7- �W��{��q��2�i�S��������2�c�[=�d��M<I�U<^����R�:&&�,��|�M��90���S`Y�x��&oԯ��p䉼���x�o��:v&�&£�䡕���DCL�B��k<��_�څ6�0�M37�*�Ʒւ�8E==�!Ϳ�F�W7���
�>ox>��I�-�'�"2�ĥ��DU&h� b�6���]���
<}�=h �y�r�%�gJ$Q�)���#<�W�X��������4�a�5`e�|�V��+�9u���Hq`�,R��1N�ɋ��[�
��R�$w��������(�"����r��Jf�f:(���@�j��Ѱ�_�`��J�؜C�s���N8�Y+����՞���W-����)���_;|�b��·o)��K�,q*��푊���6�K"���;���ՖT���lJ���g'��Ҍ��ce�:7����'���?���E�O'��}�F3h�sO.S6�ң'O޾��݆hi����w�N`} ��VբBй��WL^L��T`�b5/%�5;|`ߢy:�r�AuI��'t\X(�T=�r�T��Y��#�8���U��6���H������jlH	hAI赯w'uw,��2v�5�d�#��?�&�g8N2�Uy >�,x�/U����zx��љ�8����_����x����@y��k��*��5
�M�l+��g_��lT���D�3�;��"�gp����\Q���#��V�IiU���琍a���+�����{ͣ/s�)$����:/g&4[�6�,���?7Rg���B�ˊ�}�W4��<�~(h6����O�R�7���1��Li����>]�p�S*ԋV����v��E�uW�j��+�N$:�!��~!�� B#��5��n�v�)��ś�!dZ�@�E��s����m����-�i͟B*8��z���|r�D�U���"�K��W�2�������E���<�{��2��K�����g��MpX��끑�`��%G�J�c�,?\�Y~f?ͳ��%��^�&�H�x~f���T�3-���G?p���*T��F�&o���X�9*�#���?R����?猧�� #z����kʠP����xO�]�c��;]w�s�^=f�%�[��k���_|�\փL���<ꑮ��[��J�9��|K6���ם�qɫ��s����N@Uk�q�m�:ZB�jͯ����`�:�RVȣ�2�v��h��~�I�[��px�R�c/#|[{���������bo�o���7J��f�5Dw�MZ/��δ2�n㥱450Q�@�8�l�|��<��4:y�GSyW� �|:�i�'��I�F�r���N�p}�hݤ;%�D���Z��ɾ�_(��K���z-t�5�8F|Q %���T@�E����-a�f�\��0��}H���甧�k�B�vW�n�vT�x�l˝3�`[���� �x}-l���� z�.Z���?���'I�|P��2����8�m��(�7(���?�p��cD�k9Ew9������s��܏�V�Ƽs�nB�-#_�D��͋��:+��D�j��m3���b�)�Ѹ7�8������'�Fw޽z4��z	I�2��~{�}�w���򬚡�
(�j
��������+؆|e[E���i�卦e}�	�ߣ<��ע#�Z!��Vv�q;C��1���
si.�vfNo��Ĭ����̕����(k h*HB��7Ï7�:_�z|�y�k��d�>h��:G2�������a��[�QM��,A�2���B��*fT�t;)<ԓ9c?]E]�1pb�e�������]���bǽ0���H�I�kpܡp�:.К��[�W� EF|��Y�H�ұ�!A�X[�v1��I�J�ZCb����4�_����J ��_�iT:I���]|����M����r��Z�h�N�d=_�"��#f�Ώv[�|�{N0S�:#�?��pQ��������#sl7"�3���Jk�[��s���5J�&$��IPIk�QU�J�����/n�����|�;��0�W�%6؏6����ϴM�\���k7Ӛ��օ@�oe1��7$��_��Dn����,�����^!� ��Eq��p*W�� NJ�F<I4�4aG��3��z�b�%�'�ρd����|�H�`�����4P�����!:���˟\���(���Y}�Ht-	{k��s׷X�`�TVƞ�m�ŕSL��_�4J���-%!8�J�'��0��}q_K����L߮c��p�3\����MB�0��:��?H�T��N'�����V��EA��f�yQ2�dGKgH8M��^�^�:�#�2i�gZ͙{N�@PR6}�\�^z���!?
Hmx�T�,��a�y�r����K���"�'sN4��n�1�r{������P�;���){���`�K�%.y~�U��L>���".=���'��E����O��N�܌�J��.kAg��Ng:�az5�!�0L�B�@^�o��=e���8���
U�������>���s�7�KJW�Iy�7'���w�Y�9�U�OP��n�=G���QV U:Ф�<����nKD����&k���+j�E\�8,�e��O \���;O�3�/���[����{�E8���>��Lo���uCbּ��@�:�����t�O�� �o_U��:�B*�A��@o//����š��'��fF��J��H�){�^�4�����
4���Zf�f�ϮMa�{���q?�w���H�7}�W!�n�0e�0�����?�>?�-K��}�|L�/�l:E����E�R��|�Ex��Y�LF}7�ƥ-�%��}�u�p��L��W�b��w�9�c��d�����wsƗ����K����2P����X�Z<�JK���g>�, �|j�7�3�x[{M%���7��&��nx
���~��j0Ԯ&<�Jf?&g��}jˋ�5��o����(m���,��8C�j��:��	��dm%~Z.�K ��-��%<�*z��bŢ������Z�4��d���{��<ee���`��AL�Ӱ�~~P�ۀ�(��S�V�gZaї�*j�A�Q1$��;��W��y���߫�����h0�kk��_w%�&^��5G��m��QU�sH���1�f��U�0"�1�Y�Yh��r�f�o��DE7��O�?3�e#?�k�%K���Ց����*�[
)٬�G�(�[������V����^=j/e�X?چ;}��ٶ�q�(�e$㲧�-�	emŢ���Գp>�;t�K�
�E�,��0�`��$�vT���eC�'E�N
�!ɸ�\v���!�՝?H�?��D�j��]�]GF��`����>�h�#�M�����(,a��<��h�+�}kq>S]�w��/���� ||=me%�T�����S]�` F��SF �t iО����GR�;�ti�1��h0��gN�Қ��r�$�x#��S�ޥ�
�\�^ⶼ����b;Z�\���Ӂ}��wց����dK분yz�\���Af��18U������Sg7��i�M��W�G���r�A&_e�e&��z�%��g�+���')�3\&a4_�U�����N��o��|-�H����&K�8�"h˟ ~Ck����}_JaUo�P=���T�z��3�u:�p,���g��nՑ��xS�+��#dR��B9���#�8'�X�1 S�N9���_�k�|o ��!��!�3�[.�T�0g���d�V!��F����C,⨎SAaÍC����'ἻJ𗰰Meur�� ;o	�>��#l���P� ۰C��:��G��e�U��A�NJ����ۄb!gZ����N�Gq,�޳�WQ���<}�Q��5��Yl�[�b�9�"���+���ʩ#�Ȣ�$rs�t����
*�~�X���LvV�iw��J����H��N���v4���Ek�����
���XWvlU�XI<2���)"g���=���Q�D��>1��fT�:N�#���#̏�G���tA�����VIs�l�Z�/�ȴs���b�kv$�{&��lQv�¯{B�YEF�k�ā�z�|в��(���M��>d�T���M���j�^����@�Է4W�����u��6'L1��u��H�Ϻ7KEDv�؁adI��v�ꪵ�@mn��ճ��o(�¢���|I� h����`5�a!4$�Vf0�"��2.���Bk��*9w&F��b��	x���4N��QW��[�9���p�M�2J�Ʋ��T��R/���<ܐ��<�ߤʑN�.h�
:�a[��5�(ӕSB�"o�T4[!$�k[��F�
w۠���j��K����&�NkX���T~�*=ؠ���y{#+����3e3�:�����[�Q'��O �|!��V�3��٣"6�F��c>sÚX3��]о��93켡
�(ݗ��@E�R���>�������F
�2jlL���{��[HV%�>'��/����ๆDb�uG5F�zzz�[n�˚Q�*��4{ph��eTS��e+J�h@(�_;Y[��|���`��g�j�L��%�����r�V��GՓ�����9z@�q^-E�Ib3iR�#J�^鿿;��~I����UoJ�TX-�2����������1�e������>����6Ͽ��T��m�|�7I�b�q�_���A�(!���p�m<�x� O�!_I�\������߳�9��X���$��a�ai�J�q�F4�%����uز�������Y�<F_�3���Z5t톖���9�Ԅ���� ���_���Z�"�\(������u��4T�H	_?�m��=���B��?��ǝ���
!�̀��'	����%n8�������nV��r���7��y�`J���"�'|�A�(5RքE�8�U_ų�a��Z �����יⱵF�F�b��a��pK6]ƔvĬ�Z[?N�/�΄�����g��.i�ƪ.ܙM.�^Ϫ>\��ǉ�A���ET�ݞ��z�t/������4��ȂDd*��Zq�ł��gq��{�Ʌ�I8��k_���'AMT��ê&�[迩�Ep��R|]ztUcS��u�7�Pԃ�5�/�6� U�k�`���E��`/_�qg������s�EZ�gRc�T��lX�!L��O��Z/a/dé��.p5�+��t�ݤ��;uX+����%o���]�S��4��ë��Ԭ�=�ND��iO���ZTӲ���+鉎�.���A� ��x��>�)�������
�������h�ȥ�/�~$�]��:�0)�2׊x�
���s��"�k���^r��F ��:��
`�ѧ�x�M���_��X�"���F�{�\�$d��b�%6�]���M,sf���g�N9���f!Q�Jګ�=��f�������W�J��g��&=}?�/9:�E#����ҹ��;�a��d���(��̱:g,�	͊��z������6�(e_��1��;,�=�N�<<9�Z��e�[�Σ��nu`��H��*\*է�̧S�L`	uᅌY5���e�d2]]���^����j���4��c,l��VwH+g�uxc��W�I��.��_ӗ��dK(%4�/��bmU����c`�ڭ���E�=|k�Mʥ��dM���$-�����D6ܭ7;"*H��J�J���uD�b�O�8�p�_3�*�d�L<��(2��&��.�hl�L)�sb_�&�e3��ߐ�θ�I.9d
gT5���"$�=�����~N��0æ�[	�����ݫ�R�е�'�\��ʶ�7k;�����Bw�^���2ny��7�4@�>��%i�����M9�~�N�'�\S�%���) cK���:��ڒ����r�ڊ3q�*G�;�<�Ov�?�� k*�%&{�L�@ �褏4.���;�&�n�f��Z3�����~%����I�n��ȂP`�Z�,"��4��6)Xӣ{N�x�-1)#�<ҭL*.��Go*��� �n���С���iu�k�.i {^w���̊[�_��|��/�'�(�:��_ٽ��?�z*Py���-�^����sD\R�N<���ѥ�0�>:H��t��ieB�r��]&P�	Y^N�G\�	S��u6>׏�`;l6ٶ�!��oX6���p��"���R�4c�R�@v=B�|��l]�o0��t�Ӛ�h�uk�U�Lx<g�Ĭ��~��n�����S?�Ye�S��U�x"�$���ՎGk����#����4���������2eWq��͋�"��{<̈́f�6~U-x�GKxm�{#T�D&�*p�_���j�M���~�����`︯��|��/�/�$����v��*�]���%����KK�4N=Ԏ�>��
������~���!�7H]�6s����v)E<��c�}�j�c�)&f�c��ݥ�P8C裁�{��#:����> 6�=��}��[�M���}2c��#8ٮh����Hn�J���(R�9�x�~���x&�s-�YO�,*׫�~�2�U�M�=>�jt�[B��;BrУ��U�T�w�����U�fC1��P�h�X�<��Q��Д-wg�ɩ^�"��(�+�����yG`t��㉯����A��h��m[�a̖���{3�`�@�3)��q�D<.{����+�`�������}T�dI6s�ؒ� ʪa ��n�t�0�Og�>}���@"�`H �ȓZw�����W.��'ߥ���rv��?��;�����Uf63~{�Ũ�Հ�
�lUM��D����QQ`���5g�P�@3����7AUe�^�χz�-9��,�n��	�z�=mG�)��%0G}q��f!��)�{m
G�m5L�}X����$ �r��5%�����~-�Rm�A|Ch�S��Yյ����I��J*��CC��tQ5G� Lw<�����&��/�hǒ׌�GH�z���Wz�m�"���o٦�ni-�++����q�� �T��z��jM�tN-��u_�u��6qA�H=��O��'��R�d�S�aT��oC����w)�������_��c�l���L{�P�0GS�A��'����R?VLa#��>ܟ=�U�g*M�Y�*/+�XT_�'kog�l'R�b�{��������RV7C�I{�%�L�<K#�%�Y�'��>8dr!���K������
�D/�:�R��m��
o���g���SS'hm��%�T"���'����]���c��Hyƣ/ޡ��2���@5���������4]��n�����4��I���W�� ��z�n�����E����м�^ A�4��,��I���%|�C�[c�@i+X�#�Z{�×x靿Msx6�A����0�fq�ae3�0����>��/�� �;���c �'#2u� c�L-t5.��	7�?�'���L��
�@-e�s�S����2���|Mv��ɂ��)�2jt(��ߌ
�G�~ů�̐H��`u#g�b��[�Bn��P��p�D8W(�ɮ�%�֨�
K�D�瓇�KX����O/���������~�e�Q]�$%�Ӥ�?��.hQO#(�>w�D#DhB-��es����Uw�1Λ��V�v���LWTr�����*W�����XX�I�N��8a�r����Vr>/��2�T���No��
���P���D/����y��.�,�Л�����({������L��=)��dO'o��w���C�rEd�>Z�= ���%�7�6v00�u�;
&� ��l>��VTtcڞ�fi]�	����0�]�@h%uu�k&e�wܪ��4��z2�V4+�o� N�u"��ǋtS�R��	�t�	��-F�?�P
L�N��T����B/3MGx�
e����hQ�es�TL�1T�K��1��R���7�Gy�����I�}���eD����4���:*!��Я���?<v���ІR�~>/L�҄,��{��sDL&�@�}�c��޸{���V��1�j~��:�b��+%Jq�p�X������$�	��2a��ރ�	�.9��v��.��2HceEWB�@#��̯F�5z�}*�m�5�l#J�H��L�wV�#��R��<���F\�i���;��?CP�.��N�h�LU����#�!�٣\4CZ�E�e��� �_b3����1t�N>5{`��g�0�����l��.�5*�]�4��/���H�ѓL��U�
o���1�RC���&�EaZ`m�^)J���X�A��~��u�����.�Sv^�qR�=���J�g�* (�o�\f�#��OAl�ʹ����3�J�HM(����f#%}�'zW��MC(r�������# �[-O��x|+�0�v����Y�Ö�;�0,f��va�0��,�T����UK帉�͓d��PK�y�{1�[����,u?��+�//�8��2��Ǧ�~�zw����5�AX.U�A2$�,��g	������NM���@O���v%�l��]��Y�(��28>j��]&%$��_�pYPߵ^d���RȚ��k���Ϊ�XIJ�x�A6�o@������C�	,�B���~�b����0tm�g\7��ٶ�=�w�H�:͎��[fu�D�.��}��hO��h����=	�Ų�_�<����s,Xc�1�B�]���Cn�
֘B�<�`g�uFJ��U^�|f=�ۗ�z/�F(���̉(��ay��>[�+����=@N��J0ܔ'��VQ>��;�@Er:ؿ����ƻ�=��9T1��ҵ�P�b���������u�I��WƢ����
�EC����pc�4J
R�:��Q;Q�n��(�[��=9"�I���;Z��0��d�U]Q~���bւ��Ӷ@c;u-̚.�9�|��*ۑ@����y!��@+��D&aG�<@w&����#�{��g4jq������[;[
��l�L�{����^�������$��K��I�#�_�;H�.=�W{���2�lK�
[x:�b�q�Mv�j����k��^�ϐ�h1�����V������ ;�����rddEH����G�-��sP����0:��/��'����p�g�Y<�I���!P��MPXɯ��/�%Y�?F+�6�W(�>.����^*K��U��C�K�y����@a_!EҒv2	1.*0�L0-�]�q��:]�	�J��S��=����	"F })�\e�s�.�#O�+�;3�N���m��k���vp7h��6�y<&J�� r��`>)3�h����/�Q�kz�T>�FR ��$�kE��S㮲E0�O�dйym=��#�ӎ���� ��#8l�O�蹿�U˓�kG�;I~T�_cH�@��hڮڐ��ʉY��sp�	�{���%��u�{��) 	��w���^͍��ǉ����I��Y�o���8�-�Qؚ�����^Ti�:w�^$���Ɨ?���zS�$N<�ka�0bf	��ʐ�'សk��d���jD�����X؀@ӟ��	�����X��t4L�M�;u�<;�u�-��^V��D/� Ǯ������(��t�&+��8!C7�y��C1���U|N��{�=��(zR\���i�h�����J�pT��Og7@�g��6ϊ�#+���&]+��X��?���Hw�6�L�g����8�����e`��͔W��1P1u�0�&Y2&�g�O^r��:N/o��3�>�x�	뙉�^>Y
��Te. 񭕎�N�X�ކmS��D�9 KZ��d��<��t�����F�R|ϑ�-1�2��w �"����ht�p9Y��x��-���0);��έ�[������_T�ӷ5���u�'q�5ќ��k-4\ЩF2�9	�:^S=�YJ'��ʔ��Lͣ`��+��ey��"Nsa�L����%�@�]��e�
�`Ԓ���Ү��S�H��嬻ZU3�)Wǿ[�|bߨ!W�p���tD�����cɋ���
,��3�#2�Is:����GI���I�<���D,��a���모��}A�cW~�ԸjP(�0�y�/ יx>@)9ɕ9��|0��{Z�"��t#|�q7�����!�{g��;}f�t��Y�6�˫����g��;����Qi	�[f��[�7>(ް��]7��N��q	�s�Q�-���h,�A���ػ�k)S����x3���~�|��n��|��8���],��L��~ ǵq���2٧s����ľ�Bɱ�u�s�!/���q���/~��:���΁.�[bp�'*֔�
}����@hv��TFA(U��K�1ܢ�F`�#�8�ɗ��\~�+�i���}{����i�hK�`�R��:����pwE��NEj�X�'�RO+d�F�t��VWӍ����	�c�U�.�����B���C����.�0��| dz��s�n7�C�Y��(��e>�T���C<�b����nLa���+ Bed�H�R�2���nJ�&,CK��i�f��At�W=���p@�	Yp�lZB���|0g5YM��h`�-0����X�3s�RpJT�����Ц?�R�w5:�-���)���E>�1�-p��V2.�����ȉ��!�|k!*g�r/���3�Wzp/*�a�q�:�N��[�+���j��_���/����I���D�[c�V���Ҿ��Mg
3�d{�t�t�$��F��I��6	#����{�	���j/�>��N_g��í�����j����p�����?P��;�7��%P:�1�`���ʗf_��h��)��һH�Q](��Sx�b���n-�6jw]D0�܏f���
����"tF4m��v����\]��^a�u����bpCU�;��^Y�#�b�G����W��S`����{����4�s
��'�>C'
=t�[؃ʷ���k��XנZ��L���#-��F<ZǾ\���%6��~oa����˥�P01�2,6*��)��BZo����Usb&�k�,�k(/K�:O)�l��ޘ��G�(:����?~�)/�1��,�'�G*�/{�r�����灥���-;q>�m���lg�w���{;�s����0��`@6΁��K�>E9��������L��.,d�bM2n�kM�hK��7?G�/&Z)8�P��WҖ��v7�:������G!�[��Na�"�;U�3�NF�Q��D��B�>c	.���_@'�o"��A��ȃ� �#=��,=/>���|��QN_n��Q��ZyƸK(\�=�3g�J�v�&���^)֥u��V
�gl7yy�Mؽ?�]�Z������&{L����Ƽ_1�s�~Y���/��Ke��{�h1��ב[����r	�N�>3�ߩ��~# �C0p���Ͼt��e�ܪZ���!�QOFi�aP�0�����5*i�����|IZB��j�fP����T�q���v����P��W��������3$} g�^���8��� ��.f���}�o�2"�Ήo��S0)�=,�;�V
π�I��Th�N�?���W��=	I�0�1�-~r�렵�����5�*�b����]��6��"}I'�����I��������.9d�V:u��wϤq����&��%D�'¡  J0���@�m[3�Ȕ*6��|�Z��qAŷNA��2ˢzb+�)%e��}W������`R�ȿ�(uǔ8��H�P=FHO��Z	.>o�*��R#��X��?�.spC�,ܶ���hހbH̔�s��s���P^�� �f'Nw�+aTtC�ٍ��3�9)I�l%���kL���`��f@����G�@�Pc+�Z��|A�f�K�Z0�y�5Tz�ZsB@�
���OW�7@���έ�����L��jc"���������/�9tZ\i��#]nh:�\>�斪��8��ω�z�W���Y���x9����e+6cT�H��	����e�fuW�Z�p��\��T4x�V�G�F�Q�fd\bU#�,>q t�g4<z��Ծ�\���`�Փ��:�ے���&A�*��:&%��{ɒ��m4�G*Dp������2�^�A;�8,!J\̦H�����`��/����-�;�EՉ58�u�H���/x�z�Sx%�TLn蚳9a�[������J�Xb@>�[U�CW����(t���=��'Q_�W��=���]$d��ֱ���Iҭ��oA�(�/��X�[\|��%���a�>���. L=�$���Ƅ_\��W�9gx�E���СZ�U�*^0�ˣ3�#��B�X�GpB���`�=Q����!�B�C؃#�y�Hk:m�E�n}�{���H�����t�pX�f'C�i.���P���gMˁ��(�C<#ڟkd�q�X�+�x�����8��1�|F��S����s�R�2M勦E�&ۨ�Q R�8�D�����
���Ծ��h�����M�Ӆ�8�p�M:
�Y^�JȢs�[�~.�5��#K���><��4�!��A��$�y��$��&�=���p/ˇ=�˜�� ��x���U�Ҍ.�ô����K�KϾF��6���&"9.