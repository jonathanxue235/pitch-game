��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V����hN=��a���)�硹<H��׮��`̼��D�g�;�mR�#rj��S��k@'�q�/�ha��pc�R�(��g�F�ו�����`d%D��G�qK�DW�+X���iv�O�O����9�t�0���`�<�F�2MGJ�g_Ю3����Na/��4-^}��ru1������>�9��& c�dN���(�lE#2���Ƣ��[z��p	��lQ1�	�j�5�c���?t@W�O�`"��X\�4|��o�o�L��4������HÕ+҆���y� �*��6��.�T\)�S�!\o Xl�	=�Gar���.ū�}ߛ�fl0x��c�o$�&$ ����O�b�Q��r�)�э�L����������yx��}�JD_~.�	��-���e��>q����Pl�C?D�R��@�[m�����F�Px�Wx������ry3`�U�4&�L�0�u��]x�G=c.�8�����lm��;�����>������*��DTM��6a���:�|�Ǯu3S.���3�"�i��4���0���t�������rJ���ʚ(�a�K��"�T	7l�=C�z���Ь�f�&O�?���=�����Z1C.����J�q���J_���y�Z�#̜��X7�	!�>��iB4�ٕ��&��9=ɵ>�s>r;@d�L����-֣"k{g�c��r gq1������6����85��Ԩ��1�s��TW���t7Q�9���J�d��r��)C(�Na=����5��z)����:QuI�jց���.���Y-�bk��[}��і�̝�U��S>�j ��\��_�]m�Vd �f��KK����L�V�����dO���KS�S& �A�(s�CSQ���4�!�J�Ť΂��6Ŵu����d�`�h��H:i�ӛ�$4^*-cjj�y|�GYaZO2J�P	@,�\�;�0��2�7��q><�i�T�O6��t�'�Mf�n�oA8�-����ל�
L��_c���*�
!ri���1r�9�\j%�"����kN"I�y��k����#���L���}��3]����-�.F�4^|��>��6砨t�͛�Gr0A����#�C�[�I���T�_�+���2�@��?:���b�rb��iťW[gZdۂ��&�~���@a��<a��W�C�	c�X����3Yw�_�ڢ�;.��.$�4e��a[�.8g .�s1���=$��!�}˂?����CZ�t졁���P9Mb�9�K�Q?�7��Ύ��&��Ytw�2A���u�5�m�U�% �P7Pj��dM�����L��z
�ֳ��}4�*�'4i�ÿ}!r��?Gd,����4��3��՟�̑F��;|��k�s�r|�U�ǖ��w:�,�$[��X��X��5�@�l��X��|�,*�c�1�̈́�5����ɔȝ��$y�<���aTol�5gWZ��.�=��he��`�?7qrl�����I��y�m)k���$��G���*U�'�I�X�
���DaG�c�]v����iPo�՘hj����PV�zM1�|�W0s������&삈G2�$)0�0ɻ����կ����_lv/��+-I�����è��ALd�V'�΃aǇCk)O��B�a)�[� X��8e�X��y��x>��:���ʰ�����G�[��D�"�51@i���S/�8�����䞚����%�fu520�*�����u|�h��U�*}�:n�G��Ю*+���w��!0n�7��(���0G��(Y�V=&���r�U�qj�/������8:�%n�'��z�߿���Ln�}p�S�ᘝ�?A����}&�A���C�.3��(�#����3@1�KjqB�
�d����=\6�Zڈ�.J�n*u�,Y�B#��$�{����Q����>�k�7�HKg����?0������L�zFB@��3�%���K3s�O����%����u��JC�+�v�Ǥ�\>���;��r�`5��Bs~f�j�q/HŐ��TC�j�U�h
�<��zd�7��.%K�H��]r��c�J� �S���;o�i��j�>��3�M�Jam�-{�"�&�)`R�^cϢh��1���Z�hm!�-� gV�~�H>�K�=�ΐ۫��f\*F�+}J�[N�q�Jo+���j ukEe�/L5���w�Ԣ|�$%| �����&�w}�/������'.�P�C�̪��9K!S�.]��w�3��H�0�n��&�f�'���c��5��"�tpޑ�B�Vl	l]�=�3Mm�B��e�P�x�	�seV������jSW�~'ߏ���+���{H7�L��ئF�x���q=������!��.X��{R�����ɽ-V�v��Ʋl|�^���'��q��"���%��=buZùqݚ���hK�sW�ĥt&��;+ƥ�u�e~����Ð�e��r	*YF��
�K���QdǼ-8���꡼��I�y]9��t���U����jN�M����lo�u��樿�ៜ�Gŕ�H2'8����S�?�*���6�A���	c���6���7S�#]�8��|aA�]0%�쟬3��������N�$(a��K9���P���Ku�e��xMݽC�B��% �����p��%�i�E���}�h�J�b@�$T�>!/��9�B�1ب����y�*f5��k����8�O~���V�D���"���"Z]����u~�	�f�M����G94��dmO����8L%�������� ��I2A{$�����%T^����UӠ���5<�An�C�r��--6�=�%�}�S$��m��?��)��ȷI�
��멕i��'�=�િ�烲W��A �^�Ȩ�C_4&ɏ	���6���N����s�4~Pש'�-���V)z���ݬ&i��9_#O���d�2T��������e��ѥ��|��e7y]I��F6�gf�r�� �c�E���,��f��b�2�n�CR��t�������9����3@q@LE��'�a!�j�W�hu�kh�6b��(4IBGG����S�z,��_�#Z֥�VTv3A_p�n��G����5j��{ޚ�*��T�-_9��2�N1O�`�XrU����H�#�~�z���� 
qx�y'%��G2��2g1�]+�N"Ȳ-��f��L�A\ףU��S(;ѫ�ϑ�BÐ9���M9� ���j�W� ��{��*�*S���7���x����RR��*X(�?�l��T��B�;	R�Y֙睖�b�YCa�� �|je�+��P��Ԫ6��G���@��Q�
��\�p^�9!4�k�3� ���p*�_�xo?��ǮWT {���Ԙ�Jʈ)��������b���pA��ٔ��>��Mu���O��?��qp��^�Ƞ6ib8@���G�m����&��}"�
/'�])s�+��۪T'͔U���R؆�ʎ�ǦCR��I9�uN���F���>`H�vk����z��Q�h</�{%�8:��!|�(ųL{��h0`oo�����w���q��:[n���BC1K<��,�kY�%bke�J�;�oªɌ� �����d���	�QM1~�&��p�H�fP�t&~�2H���=:|��|f���jwt�0�.w�2>��E;�Ù�Z,5?ޅ������Z�GCR���&�r�3BT�ij^߃����&z�l�RXeYT���g��z:^M�N?��c�LO+	�Z�|9�s��kp��	7�[f�(,�I��_~�2z�����~P���RF�A#}C4�c<�fL���M6&�����)1by������u�S7�=��n
ǆ�w��2gK>'��֘n��4 �O%�K�}���ؤ�u���x/2��j�S�݋�kɊP�%���c��[�7�ݖ���!\H�O̿Y�a1�|X	$Q>Ւ�$w�ڽ�'Д��Nb�1_�"+��"vႛ���?&���"`�����K��шMgr�>�(���2�͎d��|���LM.\�(Iz��"�С�*�,��|������8��e6�a�A>�B?� N��	��/����m�����DwƠPb��JF�F���GQ���c�-[1��޼����JT�F*�k+�<ڃ����M��{�wR!!�%���)��+j�ޥʻ	�^Z�̰�'��gq'���g� ��C��/I�3�_���A�fō]V��[�Y�]�}5��_����ASjZ��ٶ�1�c��!c�F�*G��4XgY~D�v���a�{�� \�2�47}�ޣ�??pV�5�[��w2��\e��#֥�CM���f��Ǥ���y��y�b\DХ=�Xd1q7dg�_�Ρ����̨	yǯ�&TbJ��楔�[b�4, [��F}��le~%"�ӎ��#��w�޵�%��h�K�Ĵ�8N�z�(��L95w%�t��I�`��&se����yd�5Mjo���y�yQ��q$��n!Ʈ{~s�� �'Q;���O�_+���#��Dy�휨�$�/�2΃�étXV���uWf�.�)�<�?�wO" ��ɸ����{�C�l�h�n(0!>�}a��:]~MA�th��B��]C�I��2�ܪʙ�!� ~ݣϒ�r�>z�}̻��^�5�p�
7���g��T�;d%F}��#]o��XTPe`ל0�w`�}Ϛ���d�~"�Ec�_7��o`�5m��V�IOO���~iZ��I�_�"Ѻ�l,����|�?�����NZKG��sg�%sҖ�GF����wFc�H|#[?��?R{�����>Q��,[���c{9����Dr��nO�s#МL�4aj��ᒧ �M����ɯ��_	�RA\V��0���-��8G�"�_�-�qP�;������R袛G���vީ�5�~��ZW�^#���n�<���H��P�q��)�V[��3�G�*&=<���}z�!b��:�0Vq$n�R�l����+�k�>Kv�q>�K>��)G��Ә��[�=ubW�u0h��CB~��P �9�yNN,�7�KR?MZ'FY�uQF�0�ǫ�z'*�	R��Ka��9��JL%�Vg�-�h�a�Xv��-*-�M��d�?�Ȓ,�>Q,'�F]��)m[W�~
�Һû��s
�EN�ݬٻ��:~j��>&ո��y��$�A>���:�(����]��o^R:x��y��#���,��%H�RJ�a]%�}	?o�D����X�ݛR8c� �vFgw� �oC��O����uS>"�|����[�����eU�ر��ʘ�lD|�7�Rp/����8�,��4�{R�8��I�~�G MǓ�nYE��r����k���5u�t���]D^��t��Ƿ�ۿҁ��Yh-�-�`���� ����T��~��-�b�h�;\^��|�o���B�,�{�~ﺥ��V9�ob��yf��4�_Xi�yiĦ�腭���T��H�5����o��0'2�~�*���G�DT����g���?�1e+	��φ��W��M��\|Q����9�P�T5;���%�KPju֗{��!Q��'�μK�	SC���y���n�g�-���@��3��|����.�ڞχ�����=�@�;�$/Ff۞:�����o���Jf���U�A��"�p�f��L�/��1�e�HH���ї6F,z(������p�/L�ҊR�%J8sW����E�`pu�(�>�i�b���ߝR�:�����j�CHd���������*�D;@eͤ�H�`1y��3��pm��UJ�/%�;�NKP#a4|yq��L��1�t_�}��YsX��GuZ� t�a����unC;��gdi��L`(�$;p���vVk�Y �8N�ē��xe�����i\�c�x]u��1�<�8��Ibxyũ�������2�m[x��t%����5�����C&�:�My�Ѽ��(<Jh���K;{{�.Ap��N;i H�2�DL�.�jhֵ�p�E�D��0�!c������3!ء�~�Gz"������߇��4�oՈ�J��لKS�j�{6<l3Վ��_�5a��#'TK���8�������xE�|�N	���e��^��(�����j���k�4<&�pT)�%���b#$|�]N�N����.��i�nB,���;��ڥ�Rx$��οM,=`�6�m��?A��&R�WkeĜ!$
1���:t2�2t��hCx#j�rQ��+!t��Q�{�/��s䪎X��W�{�WmlF�r]�T.v��4�x�({d�pu����8C���]�I����.�'D�(덕�DO�ż!��q�x��Ҡw��
@�w�x���sc��<Tz�w����v_4u�;?� D%	*�����O�Ȣ�Ȃ� ���me�� �����箏�"W6A�9B<��4[��u*݀B�<�G�:v��2R9�E�k<�i\��s�p�^�b�BWNg�F�����	����������Y[��4:�q���v�Ǫ�|�	_�$��%"��B��uY��j����P�C��"�W9Z���$4��D���_�G^� �i:_�%������.ɤiVS���Ju�FȤ�3��`��0(�x�0&S���{�i1�Z��׹�mF3f
�s��TW��?r:is�_k�M g-�?��.ƙȍ#c�(��_K/=�'��l���Yr�K���N|#Ŵf4�s�������q��w���ϤEjm*U��T�c֒J�ߧ�Q�GdXN7�GJ%騪d��*����|�90�7l1Sq
X!p��U�C
�t��_���Q(����*�a_}[a��b;�Gdp
`�d���C8�ǔ�s ����p��p�O���F����\QG<�P

�1��H�H_\�K%�K \ʈ��;dP�v��@~��
]��QҴ�q:h.b�m���a(�$��qgִn5 �$�=��x��,�P�ҟ���s0:"�>q![�]��(v2d��,��U�Rv����YWrU��S�A�o����$��/����&�:��;��!�0։xbq��~kh��'��D-��x�l�$�w
ޫ�\�_dyy��Z�u�ؼ--��Ų ��
yU��q����kX����d�܂�?b�U=�ߜL��[v
D�Ya��R�&�fc�{�:�k�U�EYc��.�b:�8 f�f3���X�*�#���뫮-P.�V�my����߰V�Z|��d�	�pn��	����~Rj-�Z��iʜ �`,����>=ڡ�p&�_�.$�C�r��������1��9/ͨUڒ	��k��)��(�"B`�VW[���NmČ�=�pZI�0�����&d+� �i�iԬ�*bi���fDL�[���\I1�sk����CA
)�,�`�K��\�?��i8�F�8x/EȖ�&X%���;yX�i_Og����J�o� ��(�zW�s�7�|��OHɰYvI1|��%��^����7h�b��K=`o�،��ג���?;���Ɯ ��6\W���0�j���.'�$3��9��O���77-[���`�"�h�ǰ�����ڸ�V޴c��(�Iż�}��
(x��^i��D*�Q#Jzmv�R6r&gB{��=u�$jW�tC�h��[}����ɝl^o�����ú�a��d��rY	�b����*���D�J��|�󥣆r�2�Q���*(��.JЈ���B%���G�H��H�M;��?S��ChB�؏�"�֐HpƏg�v᭴���j`�ff�f���W�W���+{��H<.��kSeec� �o�TY���Q�r��'A��Y\A�b]�Q��<�����(](�Cz�ؿ�����C��hǷ(��Fw�{�6MmW_6#����je�@�T��{s�E��57i;vy/�-k�og�_,o���x["�RA��y�!;eBj�;�K/�ǥG뎠cϒyv��QP@���n��	}x[��Q�t'�bS$dND�VmT>y�*��Y��R�*	�"OB��Q{}N�-����)n��&�l�EWׅ���0���(�r� ���	Ѓc��X⇬��֖��ǖ�o��?�O��Д�k"�gh�����*��j& Ae�����:��UM)��lX���`��,b��]{Oz
~�9�[��/d/��Ol�|+UE�$`�}�=]Yv�b�b�ɺ�	q�)@�0�tĢ�k�!��=8� 	 -YK%�����3XM�F~�u6]G�TN�^�]�m�?�X�f�fgT�g�}�P4�������/���\��C�ܲ�ϐ ��+f��8�jl��(K�DQ���:-����� 9���]���T�����Qڈ>uɚ��P���D���3U(�f�O}�{�N�5/��N z�I����W9��:#�=�Sv�Q�L���Oʶh�S/�H,�ϡͻ�� `���`d˒㪩�ӤfO v1�m�{"Ҭ?�-��y8 ����!5z��d!ޯn]�5#��W��w�=���<:	ǘ1ʰ�;�^;l��1V�4+�c��%��N��x�T6����x�ԁ�=N_D�(�08L��-��%�/2��i����,��6���q��daRlca�i��
�w��ɝ��	�[��_�&Xn���6Z�{)�+p4�O���m���i����4�F�Й��{ ��J��$�*����C '?!�n�\x��_�a�о@�K�}y���P��HS1 ���J[k2
Ҏo��J0ra�%[��آ�_�����,�B��L`��/�AD51�Klk��zy�b$"����ח�3�kD=���~�"#]N~�wf�E�V���-�;��P1(���Cv�d/ƀ�ړ[P��!����8���������,(X��nܓ�%���������cB�`&AȈ������:f�?VaE�i�>U&f�rNwk)���]X��!H{�nj�C:ZƸ�Rz��]�@h�3��|�������P�>�N�e}�w��:^�@�e��
oW^NQ���<v�����2O���#�lrP��PhER��s!�{�#���6-���������}��8y��ƽ��S�m��^�E��:�'��%��JM1�P�T�����)I�f%x�(aC���Ϟ�d��Toji�o�􎦅<Yze��	�:�`.��f�B�4�;�C��;@��ɿQ F36��w65�b�n����9ה���3�M��0�[AK?�"�ԓadƕ��Y��p�$p>�5�5é����L}�⠣��*���}C
"a����z�=�;�4�sN��zM��)��r�fN�r	���L����TC�V9��'�`�n��[�r���2�(�m�O�z�E,��c��)P���}�3�%���m>�ka4�6W��A_�v�� .�T�?ғ+�kɋI�g�٩e��{�R���a����/j��hy !T���+bC�>8l�򇃽A_{1�Pf�m���3�
J��X��2w�NM����+p)��Ω�@9��}�v�j��AZI�J�����7����<@�O��2�g�Ui�Lm0�j6���^
uf�Ҩ4;�j��؉؎P�|�3&��~��ڹ��
��s��Q��`>��Ñ�hH����i�Ԣ���l��]12Q˰����$�d�u.�B,�X�%niF�Ba�VIu��]�d���"#��m�
z�(C�z]7c~��a��	���a��O/��R�Ɨ�%ag�9�k��:��%��i<˫:6v���41h�޶�Qӑ����8\���E�� `���یt	]c�ѝ�{�$r�;61>���ȎeJC�0(w�_&�Y�b��6��j���Íh2+��?���˙f���q��KK����@���O�=�bQt�i<��8�ч�F�oR��D�|���f�s�͹d�w���Ϳ�"���*���Y �;#����C�<��4�q���Y�Į�G����s�I.�ؕ��?1z�-��vi�]�S�bX7�W�=���;@���~a`�ޞ��FVZ�����m���T^���4<-Qd�$�~@GM�壋_}s�9���9�-7HM�Ǜ����2v4���%��p�F�x�t�S<��	���J�-L�qA�t%G'1^3�ܷ��h��$?��؁���wu�����}+�v����*�!�.8tڥ<_�m��f*�#��sI�=��CF�f���%�OS�܋%��K��}W�7S3<l|���׫P�U����'�LU��I�����9z���pK����10V���"�����K�|U`�I�x��>��6%~~	�s� ���*HVyql����.��) \`K]j�^t�j(�k8��}A�L(�J��E�ĺ��N.���.c�KLd��}Қ�*�M-r�" D�ޥ�ϴ������6/��A)HܐU�8c�
��8>\�� TdB�p�pZ�1'<���S�I	l�X�=О���_���1�E�����u�=���F7�uA>Ȭ�����7�%p�+e2Q�8WHh�����3�P�ysYM�	���:d��U1�k�g�z���e<3�����ST�>3bѴ~\\4�o��}(��20Q����[�������
��D�uA`�aK��qip0�.o����r��<�@�*m�t|�Bl_��.��ؿ =-8�G$׋ fI�*�D��{�4:�e{�E٦(M��rl�Frs�d�@^2[Ky�z~&�#>B[q��M��T��9��D	(�Z���4��������6�B��GQv���P�0Nsd��p֡������];�ţ��3ٞ,������d�
5����x)c(%��Ho��.z6S�a ?�-N�|�Q}�K�����'���n#�^��e,y{m���8:�t!w��).e�b�zJ�ц����#i���4�k�xW�V�TR�s*G��>;qo��xh+k���W���0�����K�~� x��We�,��GJ��.��S�tAP����&��HAŢ���=��M�4rY��,�ECfPT���W����t^��ҷҏ�p	��~E�i���L���]��A�X|J��j��R�_���~���3�{��HWF������ϐ*έ>�ǽ��YZ��w{>||N�)̴�z[~����=�+�hy�R���"̥L ��a��+#���ޜ7a�I�����xp��o�A�l77bm}��י6R
����FU�H��ʹлa���`M�ϧ/C�
����Ӏ#<�>b�5�"��(�yS2�N��(I_R��vVò�Z7w�}� #$�����ͪ��o=�%}����-3o�ȅ��������:�+���e��t�&�zc�v�����PIG1�"����N�f����E,j��N���c�x��]u�ӂ�Dv����G��Q�w>�����2���?I�g4/�2�Uv�3�4|ϣ��]W�2����B�9��mO�ﳞkcj����I�y���ײ�w	.a9o(���h�=�q�?���0�苧�cֲ�Ym��P�Z>v*�jA��E�dBZ6�0$pq���'8z��� �"ψK(�!�������2P��7ZN�!�|�S�4w*.&�S��Ըa����D�G門۩\�H.c�L�'ȉ^��G�F�	��T�l�I��1�q��{�i��~	��1T�Fsm΀צ7��a��bA*]ІM���֘��j�� �5Vs��#43		|Y�Gr�"�&��~#��E��	��o�����j	�d�}����XMQeWx"҇�	h�n&�g�yl�;_7�j,Ǧ#]8�Є�Wfzq�<Iq��1.DF�DpE��w!i���k�; ��y���vRCO�v{��BЪ�~
a��N!�|��T����h����w_!��I�G9�*�s�K:`��QpM����+~ �S����P;"��=�yq���qz�.�>Dww��A.)��2R��=�|WT�M�>'>)V�o�����P9=ܢG"�����sc�Ӥ0a7�e���(�A_./̸Y��O��;�i�۫��S�"��2�W�O^UZDe`o��ɑN�c7e�y�"}�b|��I��C[Ys��oh�I�w~������w^&D�S���v��rpX�Vv�߻�C^�5����~��8HI�B�|(�4���0��׭[�������Ɗ1��32� �F7V�}~��jI���uCBcD�ݭ�1��u&�f�=Ae��T�K}�z�x�������y?�l���!_�~�$�쎌n��k�w3�c%�������]I�*La{�,��s��66�%�ݶ}�̜nM���\�~u	��HRڗ6���"h9�D��*.s���'��s���_�^kaE퀘�r<��f_���9Ѡ_�S���=Бј,�(�l���9L�'l�t)ݰv��I`O"���pc
���h�4_���?R�x�Qq�d�Ҏ�����0s�Y��w݆a���G�"�/c�x���P�A������u�ځ��1�`G����/N����{���(f�ί�`��̴�P���q���)Y�զH��?U+���#+P� ^�&���}ggF����8ߞT䭌ؚ�tM�.�tQv�sQx%�����Tx�N��
P9��!�� up�8�y�����Jo�����$� TI]�a����sJ��p��X��8����Y{�����q/L5$=-��)�Z���Z�u��ʯy0�&x����� �����ԏr�.�N���}�ޚ2��w	3g�ˉ�)U�&h�~�Zւ�
P��}�)�t&(�(}��a��|#K^ܔ��$}p
��-U�~U(Fiݷ�N9��s?���m�qL��/JC�Wk��O�sA)�}v�G~	j�n-A�~�ޑ-NS!��38�� 	���hc6�P��Z�&����{RF�$�����E�-^ʓ���&���4���{���@<q$�zētn\W��RX���ɻιf�!���8:ɔb5"#&���P
H�pX8[v��g1��N��H��� 9w��	���S�3�Z8ߜ!��P��RĬ��W72>\�8K;�P��E���Ak�0Z�ߟ8�fB�����8�EK�r^���6>(C�.b���t[w�:I��e����))�z�P�T���)d,a'3���+�˦Y���L�A�/Bɍ�8�W�݄5�4�э.�:���z��S�K4U�J���4���Lk�R���
g8��.;3�uJ-�{���8�$T��%��26�}�c\(z��h.k
���)��� �b�Y[�{U�M������\J�ت�.�s�^x��P%n��l�x6�p�������6g>T���I���d�EMTĤ�,�j�D�x!����
iZ��_�a?AU
�}�T�;� ���-j��C3I`����ՠ��/\|����S{q%�/���C�]̿PU��!*�g��m�cz�؎d��p�/V��� ^D��l�B3�S	^�)�d��	�Z^m�������H��� �ơ��	(@�����3R<'?���ׄ�O�{����"���m�i�]�]|�\�RL2-6��+�'�{�`;��k.����U��L�6�*q�:�ZM+��B�/��ʦ̕r����8uL��ՁH�B�8���*����ǵ��V�-23W�2ᗀ�Z�4�w�n�$�̎�qF�2�RPGTm5Z��;��	�p�i�)3c�b�M�.2Bèȷ�"<�@�E���79��'i���K������+�?�f݄筮�:��-���� ���Ğ��ON��񰾶��j�YM�mg�gR��	�qq�^���4`��.�VIx;<���XnhT����/p�������~������u$K�G�b�(ߏ?=^;� 2����ǿq��5���Fr��Z��H?�jc�R�ʎ�f���/%Cf�	Ai��ɤ� �΂�
2��}�5��^��:��b���W�W�<�M��Vz�'�U��X�}�&�5�	�rw6���W������70�
B8��1Ey���O�fy��
/������dͤNX�>z_f��=MY���	<TC5�-{�ќz^��"|> �X2VA6{s��_�d
�4�ٖ�X�6����.9��b�ɑ�If�?/�z���dt6nt���.����Q�>PI���$��I��yB�۵�DŖ��.�J�/��ܹ��H(����"�!��-����%O$�f�\�����V��{�/G'������ڴw�{�09u�-
��s�?�ZM���h�!6`�L�oV27�d�e,N{g����=��)�{�X�`m)���fVv��Z���Ց/���⧥LE�F�0�i��Ŷ�:Y�O�k^`^�6=U��a���#Hq�H3�m�6@S�܂�W�H{��=��I6�>(�p&���u���a�� r��uZ���o�[MМ�Rí�W��	�:s��a�����xpS���ђ��\��@�#����c0�o	�'�4��.!k�.͹�p�e�w��_.��S40g��A>z�h5~E�`�nfϴ��K%��M��3��D2�C�d7���c6�
��@Z7P7&*�9��V�ۂ��r9�*�Ț��v8����}��w�&7YRY�+��N!枣H�]������C���ܸ1.��o.)��NS���{�̲�"��3����d[qEfle]�-�7 �<������=���4^n���[!�A2F��^�V�萲��a�dY8�#}���Ga�!&��q���dع���r�[�nT��o{WcoF��A$�;ZH;�ܨB��jy�4��5X������RZ|H�|ts˦Q� n��|����\����>��u�>\<��8��W���y,+�r��u����ˠ��&���}��D�sC\��9�h情���@[PO�9 �������RٓM)$�xA�����-�(F�Go�`./��D�X��+�w�9dX1�6|f�����d�H�FxsM6�fIJ9d���//,�"/�qcMY�k��y����X��>Ȕ�L�a���>y�]��A�hT���Z�]B�!=La�g�2�:r� ��I;�,�b�|A�*%8a�����]�z:S�;1Ǜƶ��f�leij^1:Kj>A��i#��Zk
�'�P	�ů��Jx 5�9�$�oo�#֖M�W�?���g��%(�[���)�b�H���ytz�D��K����E����}^)��v�ѻ���X�<S�����
��Zd�?�X�T@��p��Z+\����U��<���^�-���:_p������a����~���ge�mlC�{��=i�sK{�lv�B�
�
p3l���'5�V��#�^Mf�W��Մ����I�q,'Mx�'k.�԰�L��=^�h{����v�9g�(���z���3J8YUۅ`ژ�o�Ш��!�-m����3Raih����NdO����ߡ+VC�ai�< �����4�@W���v=�"���z�L�T��0���KG��	4�J��|����X����}�ơڠᒞa=�
Ҡ�BJ��O���(<#@�-DġU"�m�'F�Ho�}4��.A1r:R+;���{������pW�H�'�0m��Gd����n�?�ݖ����`�^q>�����*�+����잆Ry�6�ND��V� ��;��^����XO�u�f��Z���%\]�S�F�NHs�RP j
0������^H'���S4yxW��
���È.ߐQT@>OJ���۽2!�<}�]��[�`mY�ػ�!��#�G��hp;G����}���;��;���o����-�:,Ǔ��C1����< �O�cë5}ji��2�-���b+�h�Ա�����l���&�w|�+"��?�������]���������I�d���~���ͺ���d��|-�O}���i:u��T�f�n*O���is��TY�~t�+n̞c���N{0��.��"�Jd�~�qo���ϐ؀��?oYaE�ɓ��yX@�4�1�Lo4�H"���/S�[�I�'���WN"i�Oq�m!��я����WyO�J*([)[zW�9W�R8R�)f�mq���go�,����l��g���ؤo@�q�k��0��'�1��zn#s�3�%�ﰻ^�\�B����ڿ�L����-�Î��oqO�}[O.��3�]�9��`hԼ�9�fTs����vMÿE6(��g�)�r��w;��lv`��Q�ox�{j�J����;��+�}�T��+H~�^��B�֜���.-�룻�,?��,�˚���:�3����1����4����o�Ϟ��N�g�ѧ-�h��8Niv��ƹ7��&1׭��ǿ�F�^;ޛ��7����&��lz�pF���z�i�����T�`�De0[�\��fa�O�͜�\n�}�k{z��"D��K�VE�#�T������	0�^܋7��h��H�}�w睆!�[M������T�z�@�L���� �����P�	a��5o���l�u���x{�꡽�b��1�`N6Y%\_|���p5�
? u���u��	g�>�l���܁�L�S��s����*����\ n��5��v��g�i�3�������!��#�id��9��H�t�:���{?H�
˜,��#_)&ϓq��;K
��J6O���i���9�4�ӷ�!=l2���6�
�~? �A���2�؞�P��^6;x~�dr���cNP��%ܒ��1ֈ�9��h䵢��s?���n"N7�d�)��ʾ��eȶ"R��ɐ��E�$����������nB�~���Mt�&[D�K�M��՘�KM̜F�j%�� �l��.��g9�gWY�~l��CT��5<�r8c�?ڒ��q�,�SC�I�c�Wv����G�VA)�A��7(��Þ��<{k�y�H>���2Sv��C��C����I��XO�3�(���V���a�4��̩9s���Q�S<uJ�+3��F��WT�e�:>��9{*yt&��J~�����z�PQDK �è��-�pր�.�YOZ����`��=��ڔA ˻�Wt��rt4�pܮ��	�y���yru�1�iɢ�C�@����UR�����?�:k\c+��� ��?����!�T�lYyr��Z����(y>*���a�nA�e��-�������<򟰥չ-��������M�^�hT�e��Ŏ�mR���li�����x�˄�J
đQ�D~s���Zw�y�@���G�����(��V�l̯��X���ս;��L$~8J���Ֆ3��F������ 1?^���1Pap�����#�@����9��bnjx}D�@����w�m� ��r���R��j�$�y*`�/HTX��`���9��s�����V	�a�$����@ ��_&[j�'�s�{H&Wu�������+���;�̭2��Vi����4�o_%?�4m#�	��ߌ���eg#�����P��';p��"�ڰ�C�e|�U=R�)`��ZI��B���KCj'VN���Ɨ��H�!�ePUY����m�& l��s�{`�P"hn����f������me�"�d���kԁþr���T�d7b���t�K�V�7�>4��Ox�.�Ç.6Ѩ5�ƺ��8�0mŽʍS�|���P?>��Sdn6��'�fv��(Q
� �����Ƿ�\��W�8�7+�`�X��o�e�G�����.����*'oe�!�-a�-HRE
��o;4/i���a����;KgL���e��7�_�cM �C�=�Փz dE��oY���S�;���~�'2�=�K|2!�Y�ǊN�X���? z�?:�d�ߧ���	T�U��'�2&Z���ޢ��F�M�ñ��``�`)av�I%�?<���笇	�f���߭9����|��<��T9Ŧ)��(8u����(|�O��:Ӛ3<	��N9�A��&bg�����=i`���V���O�yGw0 @��Ab �3��F��E���Cy���z�%��לr\tכE��EO��F�6]���<_���F�ܩ�:3^yj�3:�\gۈ�����F>�s9����J�ɔ���$�FOAq��g�����E�A����'��2`=�߼/�>؁�^��$]W9$��),G�-��JBT���iߙ��Ys ��Dvu�0�o�͸�`�3�m��9A��:J����j�^������9��c���.����)�ay+@)3:�����Ew���KN��J~]�6P�mPi-镰y7��ō��7x��N���3�	w8�]���"�mg$!�<�~�[�U'j�;���;QZ\4=(kN�L��	���=2I����˵�$�M[GۈF�pq�C��:��/Nm�X(]Zy��z$��ϲ!Bv�F�r�)�6Cl��;�ؤ�ǭDHh�~��f����Y@m��R����Y�\�������t���A�Gs}��p	��;�_ů�}�m�h^KN��_�LN|��Qȇ�*6�%���	F��(��􎁤���␉��A-0��Pi�]��G�6����hn$���-]��T)�@�6�W�3J�p�D���N���?S��2�%M���t:�ˈ+�z@xX�J�)'4�0��ᨀz=��4�T�m#�pQ�JC�Y]�s���p�v_��0�끹w�4�2V$�e�c�$�}M2.�u�d��3>�W�2)�"AxF-GTN~._`����߸蚳7���AJsxQW���z�`�`�p�FE�ʼ102�5<[������[�?�nc/�e%r��z,qbw*g�A����<v#P��z-�h�f:��8��G�>�̬��y�5�����U{}Eakm�b���4��E�?O4G=찫���=�3�,aݶy-�Ӎ���#�d}���$��cT���	Jb�q��K�+���j2:C�;� s1����w��K[U�\���o�H[��
�oTesg]��^�G���j(��N�|y?�?s��Bv�PT��_*���  ��N�N�;l,��I��Y��=�#B�ߢ$��&��[�%��k��� R�%�7c5{��bգD|�P}o��U�>)�!J������N��a���	�V�U�!l�;Zs�������������j}S�ٷ2����Vn�������7� �b���j>�W�(��X�*����o�2ӽ@Q7 ��n]���v�o���j-�I;����	��s�H��)�.�)�H��V�w%��6#���BQ�&u��B04Q�2^3�����^c���d�����{l��!�~Z�]��BVM�N����F�P�g����eʦ[
U)�jVE��uܞo?�q�"��<
�����m?B�\$4���#U��l����FI�k}��3qJ���qw�'�{@����S^!��)&M�0��AD֠��g/�o�>Á��I�wyi��'���?��ZN��M��9�k@rv��|��V�Hw��\��r�*��X�Bu�z`��"%j^������X��B�j�)6�`7!|&��NLy�6V�MF�vG'@7������դ�eYW���8!��V�*�<�|޼{�H������9�D�(n3#X�{X������49{
�����kD3[�ϩ/^�����w���Y�+r�{=�.�帆Ϥ�= '�E��BuR�������î��0ח��d��g��"�?.�)3�0��>�w.�Us�]�.��W[2:h�'�����@�cu{����~]���f����#�Q�-\<�
hW2JŴ���0E��OdI�#���V�ۇBg�V�C�L*2g�p���,T'�S�;aJ;��N�glJ��6(�}x'{Z�_�P�%���{\���<����l�$h��(qU.���N�2�����5�}s��2��0L$P�U}AI�z_��v��L�	��02E��S����!�?-��������v�ˉy�V�D�Z��\�hN�K���T�m]Ņ���n�%W�L� Z����m�/1�`]1_\\�#v�0�vk�&�q�bҏ~���d+��V�'����h=���y���ul��[C�b߬�'�;]�:���L]p&Ro�炰�@r�?=亚�gs.í}pEm���TT�d���N 80�	�S�Ӎ19�jg�M�D۵�?:�x�����L=��������qc��G���R����y��d���W{�I!P(������(��8�ε�gJ��nuUɨ������͌t�I��"�+C��X�x��hs�&n�Y�\�|���dK�[�����_ξ&sҰj�9���)��t� <,a�+�������̛���}*Sa*��!�M%�>l�.�R�0��0=�q�����������_m������̅�^����M�5�?�
��n/(�,��L�Y��
v��j���l�~ |����ǧ����s
�H6��+���(���P�9ޑ���@�;�~B�6��ճ���+H_���]A��B�[��h�_����SFx'jj}�>�F5�=c{岬���4n,Xd��Qg���N/��=>�:4���t����ol�dw��C8�蝷����@F�L�v{�j�<�"x�����$F�SdY��B��i����vǈ�^LM���bʕ@w>��O����Vٱ��徤�q��p�K;�N�7�d'�3Е��e��>���W���Ip���BF�!�˦6�w��5�?#��o:�y󝁣�� ����H�h�т9.=�/(���,���)xu�B1@�e�][���k��@b��+k��m��!N�p�n)D�N_R"c��^yؽ,�~Ӭbի=`� �f�ܢ�ƹ�O�Y��O�L��eK<< ���GUkrf��e{m�A��-�$n;I2�%S6l�=�θ�U!�Ͳ��8�-�7�WW��������vp�8�u��sc��<�l+��	|ؽ�=��s� ���7᛽e��?c����?m��uxoAf���A������9[ץ��W���ꔩ�$
ב	�7��K`�N�	����E�f\���^A_��_ x��BT%�s�yÊ���BY�(�џPf�QbTDO�1�(�A��*�R8� P��o����B֕����w��Z]��%��i�dؾ�2����f���˪�n����+��C���p��I�PG�D�0����%�E1rÆ4aN��J�O-J����7`)�L�3P�?ߙ���[�j{�J���|�%s~S�*�kx ���=��R��];ې��'�ܴ�w�޺&ϖ��V�]�!��W-��y�hv����nA)M������>8:���ԅHwz�8(�B��k��|��٣����2h��_y�[������YKw������b�m����>jպ#�w�	�6hf��!a��>9�Ӿf����e�X)OB.�d\
H.La��*w���lW3X�T��z&s�%�h���S��\��J��F"Y�Le����yT��W��*A�K*�-����2U�!)��5��$dB���֫N�6�ږ����ؐg]��� K�\��.۔����"+�FBS��������ķ���d���銀ʲ�~	����@�