��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V��wg��+��1�0��"װ��_�����/$j\�4�eWL}�:�Ԕ��P���	Ȉ�P.#�/;�b����j;li��(�(�^n� ��q&�w����+�a���\��J ?#�r�xtܩ��3�}F(P��G�2�H�r5�$�2FQK��@���I\�������ސ͇�,�-�'"U��b�'�(	�s����C-dO#[H��.�N��|�9�>���sĐn��K�A��?N�������Y�j��3�0�!��߽�p�a�7��D�a��Q*c�B�(Ӣ�K҈�7��wB[�U������Gz���\\I�Fܩl�0R�T��-c�
�A+�K��j��FD�E�82ǣ��}�a��IM����lZH�am���׹�D룺�Q�9�6�g�(�p/}J���y�eV�u���\1<˛ʤB�+[v\a��t�_�Wե��g^cu�����R0D�R۽���6�D0R#4`�����_���8�٤(ߟe@�b��K��o~�t*�0H���7�ġ��9-D�e����3#�'��?�����'9a�'<����R8t6�U�}�:{�s�� ��p�[�n@�(^���s��|hr�&�kv�Jv�h#
+u� �d�>\�
U#�H�c�3c/�����^c��kO���􋁹�O=��6fw9���X�ˀ���3F����尗Ư�]\�$7�K��$WR����'�8D`t-�C�*)C� <��x̫,��_�
�9��Шq��qA�
R�eS����S�[װ�ɍ��Jm�|����y��ŕ��$�C�o��z�����?��(���K��+�!Y4o. ᳓g6uM�l��`���Dl.�����!�6����[�S��q�CY��
�g�q�5Y���C�i�ŷ�르��9��4^K=��C�r����b�+и����R.�.r��E9���8�l�e���8~�rQ\dRnK��?�J�͗�ɛ�o��V`dd�i	�WA�g �C0Y���N�݂�f.��3�EJ��=c���-R�B��αjt��>����#QE��[@�p�����g�|�����|(A�H.��>��X�
�ǥ�q�M��cs�xf����fr���C�X��3��Q��'G
��~l�ʐ)�C�I�Ǹ ��ى1J���E��_�yg>1U�v'�x�.{�=�ӂ���`*�=��"�#���} ���^7��^��vN�����.�&荕�
��/��G��(�y�=e��P����>Hd�|����Ԑ���;wR�Y�.d�6���b�$�ƴa�-8l��l.
{��ˎm55��Q�XeD�E]-������mp{-�?d�qQ���X(z �wcE�j����/�����go� ��h9�bO�����S�⿪��q�3[��z&c;9o�
@)nA\�B���p�gzV���ы:���Yc������};����M�a��p�`�/%��{A�'m�S1|��-�؞�J�N��0���7�J���i(O�~����u�\% �g�ϥu�r(��7<����י����5�r�� ;E.���C���CM�6R�a����~Wx�A8'�Ũ�0�j�� 5<��5D`�,���ِ����g��H�^"�hI�D��m�D��>)�K���\���@�ô���[ �&��U�X�_�~F�D�[n�{
���yo٧<�_R�e��^Q�A�=�mQ�V��<�D�l�%����g��װ���K@׋Zx�%[Ӻ5�i�������,}C46�ܑ�cp<S�1���O_�V��lYH��qw?|"��|�\-.���ygZ1�g �*�.�3U�MR%AZ�S���-���A��VE(\�#� �eBΦ�(����(���Z�";�a���Xc� I�۵G�ṳw{{K���m������y�Gn�\�D���Y�IFְ_'���¦��C���)#%!au!7�� `KS�L`\���
����r�=�����:Dl��v��$XW���e����/�aD��X�SXM&��VD<�r{d�O�=>���8���M����_�k@�m��yJN�&4T�H���_X	:\��{T��+�]ok�Q�q��4;��{(�n�����D̨(�ۮNy��W�����=��e�d�[�4�+r��ȷ�AJ8����I�!Rv9m�<��ֲ���Y劘�� 	P��$�ˆL#��(��H��?��BtZbc����7���Gf�oB��e$K�VR3��� :PR���/x(�}�2�̑���
���z���M��mZ��4'P��6͟�L��X�|�+��A��8�Fؗ���g9�0Iu�T=��ض3�h6�})���rjP6� �X��D-�,���'��>V_~I���$.�)}�q��y��D��I�Z�i`�ϰ�giE�����m�j#dʯ�O��Ff��d��=l5|ă��p�4b���/�⪛�.f���f�m9�7�P�o��l�{�}��uj8
�����w�!Gvm�?%��'/�H�̥^�R�⚮���k�y��\J���t�D��9��LIAF���d��Z�*����'|�s�g��#�	�WQp�h.�>�Z�K$#v�W�F�L�~o
�Hq�@Q�Om���cב.���I-JK��N}�����s���LAGG�A8P�h��r�-�������x�B=\��t�W������T�-�;18ف'آ{T�<��S��c�9��lz��A�d3��پe�^+1� \�aq��t�Po0�X�&�$Lg'������(��"J��)��;�Qw����1�c�&^k /	Y�mb�I ��8�,`ŵ�*A.*�֣Ѽ,ь�[��.o�޲�����Z�z�s�J3��Y?L�pZ�\�b�^���.�(�%V�!K,%�-�U�s�
p=�{Jm[� %�)Ĵ�!��~�Y�Y�Hԉ6��[�9-����_뎁�z�~g�3!?Eو`�����5Q�nQ�b��e����u�m�f~�6+�[	 �Fz�3��0�����!�!p�`�J ���>b�d����0#-<����L?o��W��C��� 6S�ٹ�#�<j!x��&�|����Xv3bw&{�]'^H|u�����L�k����K���4TK�P�&�d\�۷��s�3�a�y����`g3pv ���>��$��|��T���5ͪ� ?m��1���=��a5�������c3d�(3��p^���Q?�{h��A��ܥ�ǋ�Mа��/x�Dea�Ż�p�9$��	Ft���f����S�v>)���7I$��N3Ωi����~�1(�u�?N�� ���5P{TV��v�<`�0�ɳ��
��
~�.��V$(�z��^�QgM�A)��b��I��Qw��mzd������/<:�*睰2�C��T���sz��f���(ۜQ�n*p����o��#��*����消LB�@A���,�Kķ�<�x����qZ��V�++��a}_��ԨB{M���FDUx�Z����v�SX�S���}�����dǲ�)\�?��
'BFҷ�R1�ƜAk���4���-�@�e��ĕ$gc�J������L���Zj D��a����=��
Ɯ)v�-Y�DֵwU��f�~��O��C�S�E{#��.��u�آl��ھ�'uX��3�5/�8��Яv�JoОȴT�Ĥ�;5��֥��n���».��:ϋ@ׯ6.eO�8ʑ�b���_����T�@�(�A�r��)応l*��ii��`��GV�a���4�i��Q'�C�y�d����J_͘�=,��4�c#��wd�|�⢩&�����K�s�c����~t)�8p�e=�J�b~	��λ�"���}[�n$�����3^5��K�lZ�̕5��c� /uq��+�xKN���������;�j�_/V�/��DwЊ	�䜀ن��>�Lm�-�s*L�px�y�����2�F��4y݉3/�eccBv��X���)�E�?K���S�����`�r[�/|�ifmR��s���&��/4!:wT%�W1�',t�O?h�zz_��;Gn�5�����w����v�2�v��$�d7��������,;�nsMy��(�J�OP9��z�O���Wi��΅�?Q�7��Qx�4 !%0�2A���1o���-��~�m)Hu��}�ø����6{�����D`�cphĔ�#���7�:՘���nc��'
��,��T�p�ǹ�p��]�h�_�i����:Zt�fp���h���1w�<��5�u18��,4W��[~"3��\Y��ߡE�1Wq+	O*K����Tp�($&֦W�("	eZ�Z�K�%�%_��||���[3��@�3���8���i� �h�z� 7.<�}�6�΄�� sո�V\)�Y2�Ov�J�������̤��IfU��,3�.}ҥ����0��n@Z�:���uu���	3]
8�d��-J�%/��@m�#�	���P�Ѣ�ψ dD���JKA�:�Cvz�0�<&y`߲��We�D!(���T	8���L�"t[9T�[Q��!�̢�&GÓ��t#��NF#�,��0hO�s@��U�8��ci��3��Kg9��cm<|z�ֆ��Oq:-��I��:q"�T$����փ���V��Ż��� �|����M�L��G����|a�P�0��B�EX��>��SR6�Q����� �ӌ��B"M0j�B#a�2Z]Ю�E��WCy��������I\�	&�ř�S(���HF�#�
Wl�H�J�K�Â��^�>�9ץ]�Á�B��C�;�y�=v�_�-�-엋.s'�,�aU�����K\>6�;�5"����7_)da��w"	W/��;U%o{���I��aF��;I��g/A0o�(���ۚrOC�y��5=%��|��0����|a�";�T�O'�هO��)_d��[?4^j�����yzY����Xh���5˻8�#�Z����	������F�T1y�'�#z�����.�|�֜"�`0 Ղ ��BCQ� J/MQ��6.��Ld;�����\��N�������
�{;rG��
VR�'�&�˄�*�5��Փ�a�_��ژl;m����I|���f�l�OI;"��aCr�ۘ�Vo(ž�N���ľ�dގ c�bw�����QӸ,&=`D!�SmxTlH����d�j&�U� ���AǏ������$pԩ\nkq)$���1��aTD��n�*���(�W�Q���-����.QT��@>�$��Q�zl!�Z�3��z�4-J�Z��w��3+U_��3I���F@��i�5`���"İ'�����3<�T9~��H�p�~�e\�*M:���>g~mi`�j���=��e̇E(6�;�K� D�h-��z��>����]������3M) ܓ�LT˪%�2��2�χTK��ɍ�d�� ��]�pN��9D�N���E@�Ռ��j�6~�$�8!G/LEf�C���zj�׺"�{�"�K�g�����t�c|ܦ~_R�OK)����l��C�v���\�|��Na��r��F^.����d��� ��ZK���$~����a4HNhd9��O����V^�R��'��69U�D�vM�$܍e�J���m`���b ����g�7�.96aX��"LO��VQ���'I"�������hE�����I���B�Q�ix�5���A�ž��,��8Kh�`��"p��9�=g*Z�23�e����9u����s�0�k�2�Dy?��lm��N���|�\��
���C����i���c_.�B��� ��s|�}9��? !DB�!E�^h�uk��''��{pM���Co]Ƶ��}?��q-��ú�B� ި����t�T�R^����c���=�X��>�xަ2~| g��PKcu-d0 �H�+D�O��5���Kg�k+2[��hȼn��S�Ñ�R�ȱ񖨑hB>���P{�}��r����0b^��J �շ�f�5�� �^,R�5�}�®�����̎lt�G���F8�6Q�k�8�g�V>�G8>��5h%�'���;/9{PB8<b�Z��	� ~UM��rv���Z	~�H�Aj�r�Ƞ�q���n��<3O'ͱ+"�����	���K468e��V�t�k]��+��[�뾄�JZ�~��}[���ۭ�ߪT��|�r�/-m�zU>��	�N\�4��6��JW��.1��,���N�a�K�3�?�Xd�d�����NGVO��#���k:>�'��=�-&EbxJ���Q4���\���f���&^b���pm�βy�ާ�vSht�׸�4�"ʟ��A�(����vұ�&��Y����b��9�m�U��;�m���6"$Hl��f
D˽j�^7�	[B�7�2�J��N��T��墚�;5����7��TH��4������*���e�RE�<��1��~�}���c�l��Ua)�ދMl$KuۂT˱���d�q�d慏��ܪ�����v�������/��Ɛ��M���Ȗ[��Y�J{�T�ݩ��Y�L�,�)��wq�kb��}�0�ݬ7C��r�����M;S �	��*��q7�_��u��N9�9���i�0>Aj��b�����	�9�M�C6>��㷦:�_��ؖ(1ЇB���@s����X�YZ�4w,��kuC��[[F߁ȵr���!�u�`G�yˮ!˖5$K�T�{ƞ����)<��nt��v�$�HG�2�v�)�=�Z�咠Z���nP�^��S�(r',8�(��A�K��b�@���TO;�$+�(�y���u�#�t���|�bRб����.�M|8�B9s���8Y>�t���&�0�8��(��*C��������[����=A�����5s�����r��e�V{�_�~B�$�f�d�m��lNl������Xi�&�����@�[�:���Nf%�Ե@��0��^�ZWM4w;�d�>6�Mr]�v�u���1�cC��W@#
�!���*c+.D��N�v�X���n�4�&��K�W�e�Y�Ci��~��c�Y4��n�j�t��<"�[�&<J���4.��0���@�j�d��+x�acg=������mپ[d�'O��9*���,	e: �U;`���"|�+>���oZ���r�6��GY=��^2�]f�_LpC�P߇R<����~K�	�t52Y�6tE�+���ؕ��5�'�'[�7��f� %a-�k!#vm�2ڰh�t��z1�N��9�Ĕ"¦��ӯ�4�=R�,� ��Pt>u��B�W�_:й���Z���"s��GUV�ą1�u�����CT�>��n0��8GLŨ�jξ��ٓOJm�s��; ���]�Ό>���V����y�_(lI	,7��=�֧^�O,�����e������=	�l�V��-�&�ha��îqB����>�p�ÿY�� �!h��y���v�/Zf��E�'mh9�eQITIu��E:�)So4��
3W5���t��օ�5������V`��#����z\�W�L��]Vx<uk������D?�uF��8s���H�zRu<�/�ǎh��#������w����+(1p��#�<��Å��0�xȷ�9����y�	n�*�w�W�I�'������B^w]4�\k9�c��!�@ ([�V�L>g 1"y�TS�/j��x����o��vF-�
��Hf��Uߗ,5}	���f�s� VM���"X<���B�&�A�a�����a�Zk+�e��M�8���/*Bz�D�)�X~q3_N`������4��7��(�� �����7�h�u"
Xˌ<x�+�A�q( ��4_e>'��F���XM����f9Ó�VK}���"�=���օ��M���6�C:�9�9��Jp�f�ø�׶���>��"A�ED���I����^�RLr�I�Q�ݲ`68���.�(�A<Kߞ�����
�a�\V�"r@���fȥő����0D)��$3	�3�Q`Uі�]N�����a�Gp�|>NX�Vc��Y�Y�N��s/?oG"�ag&GP3t�(~�u���A+� J-bq}��ᒰ�Ts��jj��Q�-M�����������g�����Z�#�0o�6��5�}дE�$ph��O��B� ~��i���Z�,G()�V��t�8��k�@f�g�r���K�O�^o�h��A'9	��h�]\�g?�J�S4�+�'=��^`�iL7�.��[ݞ��9`Z�"�G^��ǐ+�+��>eǙ9�N������!w�вI��zf�")l.E<��ϱ���e2� ��@�2��2s�c��JRS9{V���#����!b쵺�;�U�̬�m�؉B`0=��A���Y��+�-Ԇ<>6����+	{u��~�Xd'ua6����[$���ϐX9)ITlO[�f���p�4.i�5+n��牣�v�0i�>�H?��ʮ8рCC_b�i��q(�z �v5 dk�G���6��ÓB!��j��h]�_vdyV{��m7����w�	A�1/Y��c�!�P**�TFvZOa�j���Mġ7�F��҂w�'d�:E�_�$��s.����hw��[�fY��	2���@fP���W��Z\�:G~Ӹ���+O�z����0��W,���7X��1�3�����0���4,7� ��ii�~bgJ���u����[j���P*�R��#D�J�Z,��f���K��u��"8Y�9���8�b0|3�<���႔�$�!u�x�@{^M�+p�� ;-K��Q��-嬍�:�A���x=+����8���S�Iv�Y��)����z�F߉��CթҺs؍�:�xx�P���� �*�B�}xUk][�M�O��爈{�\Ncn�M�d�]2��~�_��� ���?�6k[�{z��J%��;2��W� 0�[��/z^�,T0�?��UpV��B����(�HP���T2�p��]��)]��G`y�=hq�����p�~A�TO*aR��wX��a�E��Ħ>��.G��z��S|]�"� �W�R+���2ׂ?�*)�+麺��UPޭ0ʨ���q�NWf�#�g�|I)�4�Y(�-��R�$��E	�I%,0