��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V��wg��+տᕇqQR�WW~�ύ�	�#�9�Sg�GH*�cѧCς��J'N9��Y���/��X"�Iz�v�-�ޝRs#-��SO̒�Zt1�E�d���x�M�*C>dy�4up3ڋC<���K��a�͂ �gZ���Q�r�2L�%�'Ӵ�w% ��5W�i�����t�n�O0�딊�b��ָ�{9`�Μ8�*8��.;��fRP�������5���>[u&dv���b��;-/:|����H��VF�6(d��I��~3Ya�~�/���J��z<d09SUe�%��f^_��hL��_�����~�I9���9%��Tg�G���u�[��*⤘E�1�u)v0~.z<F�,.�7Xi56?;f��Z����v-11q� ����^�����Oho��ߦy?�������ńk��M�A�(��c{�C�� ��l�����i�u�ڒ�u;���\��wx}L������#���O����L��薯��)Scn.x��śy*OǞ�ǫ �h�Z��+��|=���	��qj���FF�B-�*�/��>;݃�`6΋����D5(�r�XF�"��Ҝl�j�.���ɔw��Y�Ѿ+
����.A��8�Uv�H�/
�7\��ȭ�,�S�8*�ٴ�@�O�gl[���혜��7��%t��F:�%/������w���kG�=��b:�,=���;1�F���5��f��_X.��N��>�QC	��n�>�R?�d�C}�;����D����V����E��lZVA�?����UQz���Y��8t9����G�pu~a[���o� K��j�������Y���&��D�������x?�#�-��Vׇq{�f��������b�ܙʩ�
��Z�3�%�����m[��i���=���s�C���]��*��s�F�~(�0�9%����T���6�'[s%ş��X>��"H2������>��[P�0'�Lڐ��g����J��<��8h�[�/l>�8��v�g�.��Z�G�s��T�O�������m���'�JGt����_����;��u�&U���pF��5�(�ִ,U�"1�pa�oio������{]W���T���ɟAY�2�-��*򾱗����&��W��Nz��Ǚ�2��z���s�)�Ss͛F ������&j�*w�_���R/ ��TZ;�Y4�;69-��+�	�&Ɠ�q��bT�OD]�J�	��#:9�@��R]0�$'#d%�{k af �����*����4"������1y�Mj���FGqb-�H�ѲY��,���Ь
�y��O$^��44LAddJ��R4#v��	-vpT4��d�C�y���6�������d6aX6�c��ڦ��
��?. ���d|{|o�,���?ɪ��bu��� �'W���+�qξfV<		a>�D��;Q�����o �Fi'(3?�H��q����v6u��:R`O�7�;�;τ�^=%��c5X�7+��������s�wn94HGBo�Kjk�q�'d����֯��n9�;E� ��ѝ�h|�fAV��5�ƬW/8[�{N����sC��"���v\�����H������'���}���D՛ (���D y�$�'Fh�;�=K9$]���4��c�Sm?�q��q��ި�=d�8��٧py|�H�kz�#�%]��a>8����[_wg�4�>���7?`6��o��������Ĩώ���Z_�v"����'�S#�֖��^�Pl-roW h8͢x�;K��5Ĕ?̶T�W�� �*���c�x"If�_�N0��p�?��-�l���JC�5�6�0�����w��F�l=L��$ŐM1g��3���n1�95t�"tm��l��C�H�1���)�j�wZ�.w^�����Y>�_��zJ	���6vD���w�@��#q�J�s��AB%h��faI�+^�*ؖ0}�6�]��&�tĵgg�1�ƫ픇o{a	���~ ����� �8A�R��u�S���5������d����4�\�1c�Ҹ���aZo/�4j����^�61}∤��=��zES�ϛ)+OM���31z��5ic���v�d����q#��(P%�,;i0����L7�NL�S��9�ԛ#�j`��qMPr��D�D���k��j,$u����P3v�
%��g<���#���g�6T���i�I=f ��I眸f�X��-����Sgs*���I�rh]�)��>�1�=�=6�Zy_F�?����n�c�p��/�~u]bו��o�C,	@�Y(��W�8�'�٥'�Ϩƥ#2۴�̐�KL���H�э�;��INV��n&>�08'���/7$Pڱf@�\��lJԨ���T�֍�M��2/�-�h�����8āC�Qt.qj�*��&_�Q2�]`���d� �	�-�F ��﴾�[����Mv�l�t�c��;u��Sg<��U^m�e�������$�����F��$W������rC�l�Ѝqx� W�$��w���AfP�*3L='�V�����I�}�VĠ��i�ʊ�6��m�);���!c�	g:�w2"���h�J	�b26���J����Q�`*Z�P[8�H�S&\4���U�(�
��@�$�$��PAr�[�=����F���?;3���ٽ��E���s��أ���v�,avp�0��!A�P������G�b�9� 3%,��HY
m)(J�v��\��E�}��O/�:�}�|���6�0����I5�g�����e�5����X�=w��o��??�A�H���}e����o(�d�4v�g|���R1F��|�%Q~I}�]��:_)�4��딾�D��gz��'�8|��^��yX{������<�M��j�p}�`�˦I�e.k�}I�[��0�/��;մ�C�sﻆGc��	�n-�hkr"�:+�N�?���������M7��4J�|է��&���O�S����m���������c�F�������ǹ�:�%)�]q���d/ѱ�a�W6���RĠ/T�%��*��F���#�c��X0>��RU�=�$�W���/� qE�ǫ������!!�ݤ.zLVsIm�1M8&*]���7x�P0<�{�-'�����2��/.O(�Y�c�_��Cz_��RNο~������{��K����S���ܛٲ11p�u�60��x�����QM��[c7����B��y	N�=`33=��'R8�s�aOLفH���|���q�t�� ◪Ұ�h�z�y]0_H�eh�}W�"��&�?ޟ5F�5<��՚���� �g�m�
U��߶J���:��_��GP�љ8��:kN�;�&i*��KЩTF���@���Z��8��BQ!���e��|�N��A( ,��ϩ���~l���,)�|���\z�-������~uA/��Ii>֚IР�lhI�Wnk��a��!������)����!��	s� p��,���`XH6��`�n�1��؀�';d��%�R\*,����&If2o��u�	c��隿7�Y�]�p��gyE��،��[�N#uR�&[ 
g�f;PZ�l�-�U�S����Z�}���3}���.����N���P�ԓ��_ϋ�K��0ވB啲n�o߬�GPht[�̦�}����o?
��d�Є��xo�+ 3<�V������H7�v��\Z}W��~���U���-S.��Y�S��}�{	gr��q�xu�W��7�����|&����h��嚿kM'd"+� BS7C�*�4zE�;CEr�|yn�"�\�++1s��%�p��w�㖸���2-�����ü�!Ja�h�G�䳻�eBJ��*���m���l�J�@˒ǽ�V�v��l�J���h�B�V��[
�	���0m�{�~�}IHB7��4E�盲	�Z�Q!�{N<g��̈��X��x������믇?K��;`��/����* w%��{߿X�z��jl�^��.@�yU��'`�L
mɎ��D{�[�{6yz�F'��WB�C�_9m>j�m��K�ݽW-�_��EA�o�I�jY�duK���S�b�5q���#L�S\�K���>=�,L�#���ฃӒ�M<�6K��.n�l�#��F����pa��RA�y�IF6���=ud�:�a�T}�c�����Ϛr�h�e�7�3��|����7ȉӂ�I}�Av%�Coz���������~ɨj)i�D0	x	�Z� m�ߋi}��dP%�Q�c�}�����I���8~��Ċ)K޴��[�,C����Yc'���)j��Pt�z|�3�	TuX ���~�}��_�s������U:d�b�1�Ó.�k8+�����ؚh�����x�F��~�2��]G^��-Q�V_n-�����-��+rL�i�ls[VL�n{��D*��RU�W,q��Ew����;60�|sO��z�!W�:��-'�ye�RG��(H6{u���y���.�߾�DXՠ����Ĺ0r)����p[xws(<]SD�ڨh��zeZN�~��v�(I���jh$���Vɘ��;�?kNF��P��@x����4�B��nl�z�ݱ�V������9�3��W�+X��q]W�cP���8ơN7��-�ݭ����a�e�2���W1��u�������Vj��[7Z����7K���2.�gؿ����%yf!��ر�>�^���S�,��F^���0$��/�c&��$TT�b;=H'�sE��6R�:�BkH���X��U�������|��L6N�O���6�BQ���^���2��U���a��`���D��O�)jҠvRG� �f�z�G[܄}�4��l,��a�'c�4�Ǖws�X/��\o���ѵ���꽣�h�u�$q�K����l6Y�\����M'����%�)<݉u���M�0���-���Y��n�"v���J}��ű��۞�%�u�ܥ:M�������vR���M	�g��LO1�v2Ҕ��O����Z٤MQ?��%b"������<A���U&:�˾���ޒ��{�:T�g7��/�M�M��� ��;U�3.U���/!E�L�.�4���Q����C�����8�yN�Tj4Gf���7�(Y�nJ��cnKϳT���z,�~3fC�hͥ�ΜRE)��m0
���6d���#4���#�4$9�~��jC�cT�; z����޻�����,F7�eR�h��������J,F�.���>��R#���:	ڋ�{o�;�$F{֦����O���~ͻ,1�QzɦIF��0��?�[V8�Dܾ������O*�)����W�Q�,{�Q�����_�� )p�a-��ڍ�`#�hF7��m��&�r�%�p�r�=�x���������cʘ���?�����rZ�I|$9�0��l2��B��v	l<-�']`۹y�篐P�_��{��a���e�Gn��]����I����h7�F@�����$�:! �ͫ���� ��%��ݩ��zvݮ���A$�"
n�Bа�==s񧧉�6�J@e���֖��	h'�5��@e<^���<�%A�7�e�Դ�r�d�ӥK⦿��Ed�nE��g��MX�+�d�
N�J? }9�q�!�a���D'}<�
�z��V�D��)6�^�r�3� ��SY�ʚjԇ芽��^���b�����a�m\��=��v�������_B!���0���� x�T.��*t	]6�Dq���1����);�s��4�N�������*�B�[} �<�E'��a\��ƨ��¿�s'	��R�]i�d�����*�� ��!*v�[�N��b-�հa��eT́��պT���Tq!f77�� �|�d�z�!o��)^�n���)��]"�۹�r9����h��G:1�">58��*]Bh�J�֪
 ���'5��~;��-�LYr)T���͒�rIR�b��.�M���!�Է4���stL�+F��4*�xd<�MOEth�*��/��~�o��T�knId	��ɓ�G ��>qw�+iX��e��=of?v*��cO�h���%j�yw��,8��X�j����Ѹ$ld���k��ա�q�L��<8��n2�T�'���b="s���������{R�cwMuC����ϊɈ5���T��AATwa6Fh?*wϱK��1�EPسfҔ��s'�99���&��v"�K��y4R�ll9�?��y����]=��L�#���H�g�*>�tF�c��������V؋^�[W&��1Uo�Y���UV�F'�t�Ȓ�&Bh9������͔����%�3�v��i������Y}T�d.2>�D��~*������QYw�{b'2�����Hai��yz�i)���SPU�b*]{g��Υ�ub*�3U$�j�<�<W7¼>�ۜ�@��fw�9���cU��|	��̅�F���r�gx�@ȫ��.Av%.f�ܼ������T��pn��ZS��Ȟ� �N�QA�|OPG�!��!�dyJCY�d6x��7��R[��Cm5�0�j^_M�1��r� ��r���V����e�y=���:��9/~F3um�NzZ��@�jb�X�J^G�Wo���iX{���*-`�e��C7���@��Z3w,�B>�B�pɜ&��A��y��2E�q���&A��?���nY��i��=!�x������⾴��>��Ɣ��S��/�k�o�\`(s��Q��P�H$Bsc�b�΀`� X���h��w(�Fw��}Q�di��9�ьR��r��B?�	��3_�K��x_�zƉkL��[�����w�K����K�.ܦ$}�ױJ�R0�"q
���g�~17�#%�]��8(R��ι��)�_���-�A�ݘ�6nݡ��gП�ڍ\j�����xx��C+�6S��#����� �3n���ů�".,�p�7�U��m7>Ԥ��%ѓi	|���Y�:ά������V��p.V1$���¢����s�`�d�!5���Ls��)�d�2�G�LHx�Y)�{�2��㼦9�J�?F�-�����y�k�	$�&�a�Oh��~����I�X���IUu��+�Jo�