��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V��wg��+��1�0��"װ��_�����/$j\�4�eWL}�:�Ԕ��P���	Ȉ�P.#�/;�b����j;li��(�(�^n� ��q&�w����+�a���\��J ?#�r�xtܩ��3�}F(P��G�2�H�r5�$�2FQK��@���I\�������ސ͇�,�-�'"U��b�'�(	�s����C-dO#[H��.�N��|�9�>���sĐn��K�A��?N�������Y�j��3�0�!��߽�p�a�7��D�a��Q*c�B�(Ӣ�K҈�7��wB[�U������Gz���\\I�Fܩl�0R�T��-c�
�A+�K��j��FD�E�82ǣ��}�a��IM����lZH�am���׹�D룺�Q�9�6�g�(�p/}J���y�eV�u���\1<˛ʤB�+[v\a��t�_�Wե��g^cu�����R0D�R۽���6�D0R#4`�����_���8�٤(ߟe@�b��K��o~�t*�0H���7�ġ��9-D�e����3#�'��?�����'9a�'<����R8t6�U�}�:{�s�� ��p�[�n@�(^���s��|hr�&�kv�Jv�h#
+u� �d�>\�
U#�H�c�3c/�����^c��kO���􋁹�O=��6fw9���X�ˀ���3F����尗Ư�]\�$7�K��$WR����'�8D`t-�C�*)C� <��x̫,��_�
�9��Шq��qA�
R�eOB#�U�e?�Oҹ)�U�i)��#�Ʊ���K�6�Mr�4�>����5�#D��?��Z	P5�W�8��u��L��#��.&�u�(L@K�L����zο>f8�cq���W������n�{�X��;�Kv=�"��di;�n+�Ѕ�5d�F�I���,�iB-�|��[�\��C��1�R�ܴ�Y1%��RNdN�`�4`}^X1�k�W��H�e��!�|�Ӭ���z�����yqC{�&���qf���0�0F"����J��tc=�˄���׮�)@c�}w��S��c]B��_���ݢ/��gk������41��wL��G���v���+����Ǔ#�e����at$��w�.M[�w�b�r:�3�H�i���v��o��x�o��JB������4Kҙ	zK �N��\4`Q�>��
E�g���2��b���*�+m���	#[�]$.~����W.��I��h��A�����?y$�7@XO9t�;�䤷����](����%yb;UEw�ȿjs�Y��d�P~������r�M�_�[l�^w��P���@����}� >˔@k��|����sƦj0|Ѕ��4��%5P��l�n]������H|����zn%D�o�� X��!���0F�:B9P�Z=]�N[)�hc@�ؓS,�Tp��|��e�
��v4i�]�;��k?��<Ml��c�۟
���׈`&%�Q�e_太!jz8�D��M�$a��v��:�cӟ�X�j����x�(%����wɐl$�� ��l#��A����cSD�݅�17��@�~�X+L����*�f��O6�����vNp��(�e0�M���p�Wo�EU�L�x�?؅n��#m}#���V��)�k�:�\���`ݫ
�/M�4�ۉ4ɱ��Ϫx�䵱S0�>�x��GV��Vk��hQ�6ᚣ����%����@߷��CԆ�p�~����ك���r�_�k'���ZJg��xC�Y,ɇ�K�?��{[���ͭ|_���bm�Ƿ�_�閰�|�!-l=��f#O�}p��Š(��/�ߪމ���,�ˬ���!��f'|��AQ
{��c��h�omrK�X$��X�T|*��d��'��&J~E��J>m�� he!y6o9�9i�ՠ�^���VC�١�O8�5�qןs��t>�t��Ÿ-���VE|Q�s��KXl�ɔG�������&��&v�D���pE�a���{�v83�d�z�zY�3t[�^���m��oJ�ZlO�a� a��A�i�17d�'�fs�; :��� XͲCr����S5ԓ�ޕ^y=������&޺
���$l�l�e q}�[t��/.�H�+]ye6�W�Oe	���b�����Ұ����ԏ���G�
K�����í7%wR���fR�1���&������?�5T�J�C�h��$ddޅ��qa�1D{ƍ�?�dh�!��z��k.��24	!1X��������h��M�O����l���TXܵ� �1�+�u̐wHX�vh���'�<G��:x�����u,�ŞX#}3�	��=a��VW��j����v�tS���f'{jT��u�Z`��g=e��i��H���8�|QT��.�Y��s��/�ٶ��o/�~����gТ�Xp�C����7Ϥ��[�� �M�y,�
�����%~�1,n骝��9�4=UscN�aa�d�M��r�6�*���b��{�*�)�2�kOof�,c\B"떑���/{��H��8V>Qӆ�j{�R~�9^��=Zʬe��}�^5��J��N��	�'[m�(� �&����szEۃ�^_����+��r���f;"�j)(��}?���-����g�<�ޤ��v��8�h�]�8d���&�k�@%��c�e3�}@�֫��k�܉m�ԅq�%u�C����Y1�S%.��% :�� �|�p�Z���߮?�ݫ�U洼�=D��=B��$���h�Hq�]aY@��{�DV?nIH2aYAx6�ͯ^���^���m�1z3em)cS�*����79x�?��cb�$s�Ζ���G���0������|GK�F4'x߂:>���C@<�1@s��`a�t��0�0��y�I�Z�a��*�i��b��e:��$��Wm���'�bgKƒ� &��0���L����@�u[�(n:W�,(\\�ͫ��:ӕL`�l�,ZJ���'��^8����VzT�Z�K�M��/���Ŷ;ö1c��)w'�]>�sbc͈�X�aA�����ӗ��]TM6����A"�m�`�U� �xH�'������
m�m���8uE��ZI���g�ܛR��d�-�U��,Q���`��_F^��p�o��
��(�6�NJ>�Dj�Q%�Y?A��?>��Hޫ��W'��V��`ԇ�u4��fG7��Σ�r\w���Cɴ*�˦�?���B�����|�sM���Z��3��ܩ`+���l�̪����}�#�p^|n!����C�J\wy_��"ҨQ.�nlgCqD�ڦ��ů:([�w����S�a*��I�B���6t���=n�I܊-l�P�]��*XQ�F�oP�R4��f�D�>�Z%�WQ0��6Q�.rk4�(�ǘ\KE��>ǑFpZL�{+xUZ\I�X�&AcA�g�'@A�ҤӢ�v}8)O���BL��`��{Gj<��-�-4�`D��C�J�DD��&��K��|��X�z�Z975�%QB��~^�@�Yȓv�ӭ�Yv��,��L(�NW���(%+�a���=D��蝲��s���`v�D�{�+w��n�N!��m�����c���	~LZ��1;��dy($�I�#��G��,�t')�1T'�R�<+m��~]�
��]�3#[��^7ŷ���Z� �ڧ�<}��N<i�͊z���E��A�b�.c{]��~屒�#��;�R`� $b���Xk,��Ԯ]vŗ���!�i��|�B�|]�d���^\�9b�G�,URp/[�����"p��e��c�%�Ғ����y
��y\�2�ݻd�Y�2�U�>
�&�i��&(�����E��m�'Em���V�^;��H�W�l�魯��&t����IS�x�B:��ڏ�������d!�`=��H�/�;��{��+��<����c��dp��U0��OK�z�6�F����Q��pG2Pk@������4�U�Ĳcσĉ'3�1�~�B'z�̴�_�oz��B \Se46�D��A|�6ٖ�H��������v���t'k��J�rB��}�r8j5P�E�[	�_���\�Qlꬁ
:�y&����l㴪��J�r��u�촢ҝ�?+������i&�où�2�AF���v=��rʱʅ��z�.�[5����]G�m���9 ��c3)E����M��݀ĭ����s�7�;-IhIy�t"��TȘ��E	B�~i?� �f�ݶ�L���+��x�ՙ_�"!�SeZ�Z���n��*�c��ḋ�=�'}�{�a���{ؗ��'g��i�Nig�K���f�*������8m|]�7��HM��C��h��>�#7��D� �FA��[�T��to�������V�ѫ�s�Ƒ1"1�q�|�H�*�x$M�jQNo�+:p~��S'����4X˯�YW	�a�&Ekh�i���ߖ��wa�����ȝ�Z��w7	c���	�eu�G���L��^p׮�H�h}�9*rb���ʫ�v���N��|�:p��x������L�P�/���N�MH�ة���.X���Ձ��[]���du,��t
�OB���\";Lg���]�V�(��AQsjX��*H��O���{h�����U,��=}�g�x|��>k�Eh�
;�(ր�H��"p��:0�3y��:�����.��8�o�u�Ri'�6���!9�s�c�J��'5�&�'��Bs&�B�q<J�:��]\
���3D���duY��ύ�$I��ĽP�|�ldޜ��X?&v�|&��7	�������(�;�]�ڔJC��f]G��O}�#�*�:���[����rٔp��A,~_ ��C/�Ɍ��<a��z݁|r���V������]��8��;��p���L���1L˲�y�/C�J���.#;�I�ۜ*^saF���Yhɖ��ށG�R��Iݹ@+¶Ȱ�5�&r"	h��(�9�{�m���7���1��5�T���[2@�B�:�HUhD;�6!�D��Jd�A�E樁+w�}� ;���},�o,"�v��a:�M21����'T��>s���(��K�^�p�Z��F��b�[}����\Έ�}e۶R�.eJ�dAJ4�赟\�R&S��6���ߗ�S ʋ��~����5�K��=�5��|A�d�vq��lg>¿>Ө� �����y.�)U���Jĝ̨Ma̞7��wz"����G�#��Ƒ�J]��Ӱۖ���:f7b�H��8��~w���{�C�A�m���n�v�
�7d��[9eBz����䫒]w��틩߅������RÔ�ę!%n}�����1ވ�*g�B�T��H약ks���u�솣�=�/��+q�'�f�����[/N�v�%n�1Q���ΥO���mމl{���M��W>��+_$b�w@�]�wkx"��g��c�$ �@0��a�vC%�L��p�:P�v�E�D;� �����u[4)��`��2��L��8��`�é��߱�����Bb�4���e�k���"�Q��1>Ru.�+��S`���Lc~$7L���k���Y�b�TD�<N����f�gU*H(�I��
���Z}�m�]���O�b"#�e� r˄ǅ3����_�<b�&�k^�r54�ǔ����H9-@�{�f#��t���D��V��_:w�%ѽyTzqF�P�#�bX�����"�c��� ']�"���#�kf�I7�%do�BZ��?��kor��3dԦk�n)7�jD�9<�-�+��qu�����
)�垱�THk�/�qP �z���0���>����������D��F	��HH�4�<�^5	 �D���]*�myr���-�&���޼��my?2]�C�a��p=)��`�G��g��g�m�m�i��S��{d)fN
"�s��U�D���4����R[=Qk�����{B�5�!�{w.�w� +��
V���u��R�R�A��D���H�e���<~q6f�S"�����A��a~�@@�o�W]ճ�h�K8�N�"��I��W�w��T�z�\H/"�%M�4cv����b�b�AI;�B���V���Q�[�o�<�oυ����u�l����0<m�q�w��^�Ae.V���~|�ӑ��gwp�񳇏uQ�u��&�odl�-|RtbCb�F�`�F#+<C'�eg��Qq�/myO���٢]�E��E֍�]�R�����i�t6��D�o(����+g�]�Д�x���W�v��U)���Qzʀ�:"�W��ǅd���_�e��(��Я[��9�h�8!�r�&�l1�~�H��=�p��f��Z�S�|UX����zo�i'-��PX���	_�<J'�vz߇f�k��`F�����xn�e0(P/حaa=��+��8̧��D,�*%a�D��c��q���^�2<�s&3!(���s�r��)�%��ޘ��ػT$�Hψ���a"PE,�<yB���*f6�ϸ@�Q/�a'����Y�t�y0��)�޸��'ߘÎH������OFw��Z-���	��:L"�R2�t�	#������ڲX)軷rTH+�;�nlĄ�Y� Y9�rߔ���W�I�CTѬ�8��0�)B67SEN�w��,��k�̓u�k	a*����»�Bl��ip5AD�`����E�Q.��x�D�ٞUg�7+7�W��s6�r�}X�L��a��">w��Lg�z�
��>?kv賐_mqv jFk2,V\�7$+���l[n����FŶ:�V�h�'Le܎�يg�g��h
���V����〈�W<����wd���O��V��c�g�˳2D*X?m�_�K��,���n��ݧ-{@��£ǚ:i��{ca��3���(�\������IȆ�ᒋH�x?s��Db����#��$����т�-�8��.�S/��f�s���z�<X�'�J����N��	<��� �Yh�k�>�Z���ұ&����M�P���y�����m����Hk��ە��G�'�K�.qN�$�� ]�<�M�I��MFu�>�U�&Q�H�UDXb;����oe���*���x�
=�;8���Rv0	H�l�T�����"�M#2I���<rr�X���(R46`|�UG����{��4t�5��,A���N6�x�4&�5���=ا��>�-�떡��!1���w���ώU�()%F��=�S��w%*w4�.c��!J=,������*�Jv��������+/	( ��0bj^Ö?��iƈ1ׄQx�!��hm�H~�4�J]���xX�(��������B����w�lh�űW�MF?^�.��ϻ��.,����a{9Lb$yQ�z\�ܮɝ-����=O�.�U��}�!�G������Ӻa���]^�h1'kl���/5��g�Ũ�ydry�.n��mK}w�� ]m�6yO[�$��=Q$H���j��[��RO<��7�$S� �.ŰO|�֘���+��`�^|���Ri�64��p+�,�(�KAβ �q��g�N`g)W��� X�����2Owsu��	�ۨITu���-,�:m)P˔���^n΋�'g6��
�)��hO#�ڤ�=}H�
%��7p�	.����H!�)O�ޔ
x%(��q�~�����7ͺR3�	@�H
�i�������ե�)�
o0[ F��)��$(�vzA��Pp�Ch�o6$(v:8�*����¿���X)OՊ�5���h{�n����㇪ļ�w�귉�Sg���O^	e;WfFP9e`#�'D��$����X�3K[��'T���0��0�DVG�^!ə,M!G�x��MбUh�ҩMMUt|���l����>��Bak�En��®H8S[��P1 �'�˫ѽ=i �>䠪�FT���D�c��xq�ɒts�~,J�Ȍ����DB�� �1�o+:�v�Blq����[�A�F��@��S����ϖ�K�F]c���r��G�l��$cp�ʼ釠U���Ϫ�i�Sn'�-#�����u|b�|X�(�27��I���kd��38m�$��޼��S����	�Y�� �<�C��M���i\ƹ(�|B(.���ŰD���wS��3�:QE*�ȡa8�ӱ�{��pi�5f�����h{���0�E��%�$1/׺��Q(�ӹ���p�z��X�zLeX�P�2�Û��ٻ˫��%ػ�F8��{(
#Cigj^e���h�����Z��c��3�>c+йu��u�%'1��e�*/�|v�q_�n���sj��)���M�.��M�Q�����A���s\�Ӿ}�Y9fj�lh�������z�Y��}T��w��C"w��1���zC`�����j�x���1��)�R�@ۈ1��4\�=��K��W�����Ze�wR,0�9��Sh�o5���n؊ǹ� ��
	��rF2Α**H�uq�W9��CYh~��BX)�+��-��>gNY1��=�gmm�:�D\��\3�>W�m��	,���a�TR�oa^�`ֶ>��k7�)���K��/��n]����\�����׽o���T��� B�z��9ʇăb_N��%\���t�v[eo2�����ɞ"���I2G��ۋ������;֠a����G�*��s�-��gD�cHg��qD;D��X�ΩR���غYY6�Q�H@�`�J��*�{�a7����Ꚋ�2L��*m(�$�],uMz�쿷mѶdSL����F|Hɫ�7Q4����$�j▖��,k�:�a���W��Z��[y@�������m�lR;�h�v;%�T�-�18qY���J��:�tZ��
S�����m�I��{Qm����������6|Nj�,j�R�/a��a�@�m��7�fՓd���@�
�J�<f7|	ƍ~�	�ެF��畮�g�}�x~�[-���˫o�e x����l�{b`��Gi$n�?�|����,�O
{�~����<#�{v�)y��9��^O%eJ�l���Q�	\�kľ����^���C��3 �$^�6���<2l$�!���ԉ2ݼ �n�VdJQMU�nبD.i�]Y�� E'z�?(�@)�{�8+��\w8����98�)h�����֎E�Q5�>y&�m���9����.�+��r%T���,�l��4��z�^T!��d�b!���\����g�`\tU�>����QT��n�/
Ɋ1(�)��n�[Z���V�dc�d�إ�ݏc�t�.@-:�C�|F�Mh�%C�M�/?���M� ��?k��[K�����c}�������h)$LK��w��'IW#����R%�!�4�k6-(0��i`��mʝ�m�r���ߔ���O���U�n��N豸&���,�i���@���F��,�B���r�8�1Yb}}q��m$�FJoW��t�(7_��be}ue�u�Lܡ�f���
�Ox���^�%�28h s��lT�A��A��yA�w' �sEiE�,�����k����CFS e=̜9^�eѪZe�L����1����F�ê)�J+V��gn|~X���q�%'ī��l�nD�\>�yUK���=$�Gz�(f�!p�_�Ka0�]�߹�J��5f�[y�t���O�O�'_N����$�-��L�w�~Θu]�����F��f��PkM6����R��f�0�M�W'��}
I~.}f��I����%��Ec��R�h6���5�&�������Ȍ�a{�Q%_TETF�s���<wF����Κا���������&�3�����k�mDJ	R��.}3��YPp����P�lj���j���X"��ю&��cN�����m��l�L�\��U����\�Ӿ��ۓܞ,͹U�����,G� O����'��08�Ȯa��8��e��M�7����@��� h�eM�s�Ae��|�X E�>�R{�q�y�t�>������R�˙��c�?�$=�X�Jf m��$^�I��l���3�`['�f^���97���Q�PIq�M�XB�7��u ���b��C��{Pyo7i"�ot�S���l��M�(���<���O�F��%v3N�����;��=�s;���<�+�5�WUSH���K���
(�q�Q7��~�p!<���Όn��yR�1��+I j�8-v��!ݙ�<b�g�Hϼ)����S��eP��h�~;ѓ��-G�铝��IΑ܏E�ez,�B�{s�oM��veh���.�$x����:As<3؉v���ي&fc��w�<]������K�qY�p�6~���q��q#��1��ִq&����s�/1�&M��\�kR������B�� Ϲ/W�tЌ&U�s-����&�ZA��ϲo9�4(��u>S,b���;"�[�ȃ� ���I�q��Zk<C�_uM��4�z tąV��`����� f�X힖ƾI��Zc���h�T)�R����۸���z8~�Va
TKL8����Hu��ÌB2�Yy��K9��,KAM�m<O��ͻK��З�*��UW?�ih�#�^0uz^����
JFA{��]BU*���C����"�L�T�{�mX�C#�[-#�{pa��萄�U��8�ݷt�g�P�S��u�Vt�K����!t��i��T��Q�w\��A*4��݂���bژ�sA�$�ݵ,�."��5U��P�d�1	�t[��.���ׅ��h_��qXG<�e<�ڀO�,p�2��h�_�J�opr@�ƻ��� S!U@��eɁ�1y�&E�6��u��ޗb�S�������k}����4�E*g�JY�T�0]�0? ��y��3���Q��I]`z�N�MB]�\p�ϛ%Ӯ�A��⫊xGC�c�<�n��F��4���D�=��T��k�)��6��ݞ+Y�{<2��07R@Ӊ�#1���pLd�Y��v<�����GMa5*�þ��������F�/���o�kվ��Db���ϵ�r��Cx�((��t��2����������*�|�+wb2�'�"�x�8�Wc��M"
I}�]� ����p�{��v�#`C�EF+�&�	���y��\K�<��d�F�rs�����~e0�|`�,i 9;d��6�����,��+-��wbV�)뫺����x �G�VI��<�v�B�����QG{9��H&E ڣg�-+RU��}P�0��s�C���L#q��!chC
I}�'�'�q�Lb��*��������/(��X#�~�I��C[ V&k�?�ƥ�Ŀ:Kv��I���T�9=���ނ�أ�b����w5b66�?jʂ� tjA䠝�S�����m��~�/�`^��t6k�&���'#e�Y��v��;�Ì��.�ļ�7F*�QB`C��tʳ���cL������Y�M��Aco��v��]7�ˠ���u�t�]"�*�},�-#�P�M����?X0�zcprf��L�r��&G=�Mb�]�­xn0;^!FސUz�������nͪ7��'��E���y!�\WEZjlW=���UUE̩�䓐s����q��y��w��0�T� ���O ��>�c]0t��X��'�K?���=����!~�mpM�=X�cal���fU�z*����$����5�E������lJzRcSa�r�?�~F��e�n��j�N��OU�x���v4�_K�vY���*�n<����ȅ�i���Er�Q�NN����ő�ִՑ�t
�S_�dB���k1�ӳ��d�g�uĕ�1�E�H�EoMPy��Q�o�=�f�q DȈM_�"�?C6xH�?F��l|������J�m�UɧE}8�\�@!��#=D��b#��#��C;W��_5 O�%���ǎ	i�i��ͫ�!,����45m�Z�\�ܠ,EjWK�8q*��:��;���U�D���*&.\�T�&'O4�iZ�U�3a[uIF)���s���ik���(q��U�
�fр��̐x�c�j�V)9,����$�&�洨IL�.+�s`���1P ���j�4��Uş�^�D��}��dpF�4g^�����8�xu�No7�Ԣ��7`g9Y}ZB�#�󾙠�<L�h@ #�yм�uA
����f�x��Q����<�u�|~�SbH`���7
���J�.�X���{��;tu����N�#�qΒzv�Ʋ�dhB)qp�_$:L���]��[z���1���qz�6��/�Ƀ�?�e���PC/U�����A����=��(2�/��{�q�^��¬㽧��po���^>��>��=��_͖/����n����{�7�=�������_K�.C{� �&8�G���_����	��E']�A��5�@������<�	mr?IS���{>M��pz{�ꋂ���X��G#���c�����mo�	����w����$�hxַ(Q-$��y�4^��3j��c��B ��v��o"�H��DA���5l�\�6����ϨZj�K��V�q#q͟�eW�~�c��S\��ܟ<ֿ�>jKdS��lQ��?��2�dh�٤�wX7�2���kg�����pK�=�'�]�wg�N��&R?b�����:����u�F���G�ƶ�[响��h��h��R��c;�iT�WZʋ�t�J��!�ȝ�f�uZ�ƌ�p�1�����p�v���6�rq�9�0l���>g���Wz�O�D�X��0> |�Ĝ\y��`�n�nхp��]BV�5<�I����IΆ�2�;�gn����W�2��X������銦w�L����9�0J���G-�Tl�n�fC��
e����d?{�A�U��6������V[]���w�=>�Ԃ�]��T�	�j�bv��M6���zP�MZ��!8�� ��)&���y��	�<~��hd�7-< B'ђ�|�fG_ީ���'�V�v_��$,df��8R���EB��z5���.Y��v��w���t������]-ZK1Ύ4�O :�����:NL}��D&-i�(
MKf�$���d��i+]wLNs���q>O�~.1�����d�X}#]}�g��Q�S(hB.6@W�)"2���a*�zT�`�m���E�5��0Qh���>��ȿ��d�i1z ��ۉc��:T��m������!7�MJ��0>�"�^*�v���g��\����[�"�⿬�/�[[�<r�ш���}��?Xs`���L�`}Y7qv����$����mU��Ym�e�ۨ��7T�h��l�x%��E��Ǧ��e�y���
��uK��'��U軡sj�O��'5)�k��+��T��;��Hw��	c\=��o6��z,�~!dj%<�:��^��~7����jвj#ϘѺyl����8�6t�TV|��()�[��UΨ�e�m�,��D�.$�E
(�uQ��ʭ�ʁ�Da���g�w�?ѥ�����&�PD鯑���R8Kٟ�:��p�}�ܗ���~��[������F��8k�-I�+������p�E��� ��\>x���]j�b�L�V1��IF?oJ�7��|���̺2����ة�mV��o���l���,���2�Z��˂�5�#A��,�Iᒂ�K9u��˳
�Gj�"9-���!��t�����=�L^T���k$i/t�}�xb�,�x1P��l}*��?�SJ�|Ja�ӻ~v�eQ��B;Ý��2̔i�Ħ���Q|�mH�����(��Vo�Y�L�!/���+!�_���GGz\!q�*�bW81{��"�����i?րF͵p�P*t���,R���B�q'�m) �V�%��OC�VrQ
	�����R�2��^�ӊ�v�4b�9H��NO&� �/K[��A�5Xۨ�&'��L�"&�6Dᧁ���M�,"K���  �!`��xU�:VƢ����HmRh���.u�'�,�K�pp���d�t�>��R!6,��w ��qP{j�&��-�_X'��]�m"�]����|di�����S3�z��/.�����mo�)��yC6�*K����JQ�҅|<���sݨϸ��-e��7Bes�]� �uG����>\���ph�W�'���a�{��s�B�j���C��1���F�'p#V-��Co��~�L�I��Ԓ�\�m_��ˍͧ���<� �A\͕�K_C�_��{372`��S��f�P�'��Y�~ �v�e������"�z�û��� %^^��T['��)���K/@��K��߰�%p�Dж�n�g�/��?��
A�����&���:�Ҩ���'�3�	X@  )�����$��&�Z�x���Re������!I�9Ǭڒ�+A_�P)?�1^��dQ(A�7}W9j%���99m@&K�(�"�DY3<ї����R	���q��"W^��;+W?�1�l,�O�z�љ���E����F�?�-��~k������_��־8�:������%�S��o�����);���9���֩K���_w�Ş\ǌ�(�a��DOҵ��ze�Ü��1f�=9Ap�kg���a�`Ŭ$���lt��ʈ�2�ᖨvs�Ąc.Ʈݡ`��Ys�	?}.ۀ��Y�vķ+�;�����c���r��J�����{��S�o�� ����|��ꉨ^`d>�_ܼK�D�Zh��՚y.��O�;
#n�ޞm��Seqr[���0�	�L��$�y��9L���	��	�y���=_s^o�±F���ꄟl{"��{����n�$�`�Bpj�J����x!kr��Q+:)���FQPkZ`��Q��qy>��6�CdV�0�$O3�_.��䎥�q��-]�x~
k��v��r�m?��lXU���Q*􁔫Y�q��
�w�:���?i��6�Lf����^���u��俵h�"��|B�we��BӐN/Zs����n�	��M�R���N�,��GuN*jjʧg�
�_rm����	g7x� �(�fT�K5�p��D$��3�7�j1:�<oP�Yn[���q��P|Q����5B#��v���0~��f�+VZ?���3��Q�<`��Y��6]��mx4�V�	�_���(�Y���t��p@����G;9�`���;�@!ɜxέl@muly�Ս7�j���Q����+����/�aRP�YCd��B^�0>�}P��]���‿HR("O{��!�I�d{_�II���r��¹�,���%�t�գ�^�5��]����7�֗,��1��E����9��F��|1�޴N�J�e�E�X4D�=�7����|XAW�b��Z��=��3�7{#.�&m��!�_z���5F[j�����ǔ��p��C�X�S�ܦ�R���o8*qW�u_ ��_T��T4κ��F��r!i��H;�B�g����S���2��۠� �~eF���@�kW�ZT���婘:���lː�3;��5�C?�c;3�Lw�v�r��&�l������!�͓�m�y.�8��������%������bdPYV�KIC���]�/�u|�R���!�b_�C���ي�Sza���� y��8���6�	Ю���0c^s��C!�}:�|�E[��N��?;�%��me5w13�7��^�a�-w���U_`] ���g��vhS;e�ͫ� ���S�k�e�p�D�Nͩww2U#�2��9&g�����C;�3 jJ�2/���9����!�!��ɗ��|3�G���T�� ���s3�k��ק�����Ֆe*s�;��r�he�:�*��Q��8j�+#�������u��c�g��<~X{Y8o���5�#$�
\�닼��2.�a;d�P�BK�p�ډ����wP��u�TRR8FPMb�Vl �����0v�k�1aʅ��%b<�W.�þ���k��,t;:��������Lݡ�~ǽ � ~l7�.��w��2�3
�_���|�_ H�7�G�ϴ������0
�!F},:������&ɫ]�(�R�G^p}��?Uuf��>�z�
�Oǖ1/���Z�����M*C��X�����)jL�Ŀ�V ���w��ݭ����,z͌r���0	f6~�.j��5{��]<VOx����
��$���� ��ۼ��_����������`�A�> �����N9��?����U��H�9���3"�V��ߺ�������,����9G�)�_`6M2�����#1�hIU�A��k ��Bk|S.r?��6��̓4�iZ�Ok��>���v>��������HT�H�O�JS#^���ѿI��<U2��mȔ���|���ِ$5k#U�n�Fzj�0@�l�Hgn=>❃$x��Яyǿ�;N����^	�]<*ǟZ[}�h}���0� ���88��$)��p�� N������E�0�b��W�3*���*:�`��h���c�h���:7�*�o�it�il�b�+��F�-`IC��0ne���3�X���5r�v�H�CLĒ�pGo��R3�����ĉ�}I�,�g�|�!k�������7q���݄A8���=�S�ѻa�I(�W����}͡�/No��OlL�pdg�~�90c�<js�5`,���i��8�a�m<+���rɎX�d�ZX9��T���!{*�#�Ә�*��U*������m+�A3�*�S.�]ɏ!�f�MQ��o��[�\j��au�8&`F��8�eOz��i��O��r�r�1@�A2�����Dh��[�2䎔�7U2�-�Ho!�]�+�&A�b
�`��)s�T�~��5��U�>B�o#��lL�����2�]��R�q����wB8y�;�"괺��[r�L3�t���a���i�O��ك�Rv)���g'���n���2I�S�	��!���X׵+�.S��Y�n�:=t�Y��m��x�\	ǚ1�4�e�����A8z�^N9���_'��P��(������ Yy;����}�H���|{$e�y�w��ǃj<�]������M<'�y�H]~3Ip�B@��&C�Tv$�|�@�}'t��k�.���}��r+D	;��G��ܡ�o�HB5����9�7�S�����mG��Z�L�n��O�`Q�E_�/�N7��M�����,[kI_��G��5�����e�x&��@W0<a�i#xO&�J�_����ϩ�k p�?�Vz�ǰ���?�o�w�����7�(4�E���]4�x��4n���x6��d#C�!����i�<9���z��<T��~�H|D�מ��9a3�'F�#�����3<C�Σgz	2ff��m�ul�+p�.����di� ���k�Es8j����01�é�yo�P���h'=�Q�7�AVA)�1eq]؆楚�Қ��'�<D?|��k��3f�%������{O�����3g,�'򡁀���iAs��2ƞ{�:Ό�铱�~�6�gn�+�(w�mޚ�攼��d\���BUj�q$՞�6/��1�C�`���pu�Fp[�E�K�����M�Q��n}e�I�DPB�#��r:s���)�[�\���R�+W�zҋ�����P��W�ʷ��+黧�b��S�֌��&f8g!�eY$ā��U�d��LI����Z��x�[���[��p��tZ�3���Q~-�k��^�H��'{w��T\�Qq)`��f��aF0�%%,�$�I6?e�*n�����Ԓ�cKI����(�ꦤ{>�o����g�xŹӤ�&S�5�:Rǟ�um^�dvx8H)����=�a�!����vK���j|��Ҍ	(��5�&�"���C+�/�jT�C3�ޙݭ�&�pmXw�T�݆���Yܿ��6�={2^?iү?][��kt��RND��܍'�1�9o��f�0�⨼|n��U��o&�eEK��rG��:a�����0�x�c�S�5��/�f�p�`1�IV �$?yf��i��y����<��q�΄�m8SG_����Jr!C���Q��hN�u�R�>6@4*>�y��+w����<��`{�<@�S�"f|45�C�W��߱��>`��N��­2�$*�,�M�HЎ�0��2�D���R��W�c���������1]%[��K�x8y!v�P��K8��usU�#�s��;��Da&�4��|�~�&Ƭ`��GT7Ķ\� &�RR�8�����󶢈6�"TlxJ�`��������ʭrS_��`����~y�s�����^LM���dDt��U�e�i׉�B�W��1�k�gwP.�[���"���<��$���kL���&1�p�/�$jK�f(�#Z��z蓚{�} �FAE2�Ց�&uz��LW0��]Z)}������w/{Z��L_\��2_l'�������3�Ȧ��Ǉ;��[��Nb3�rf�l�:EV&������;~�_zYZ�=h�jf��;��VN�o~��{[�s�DC���F8�;� �Z���|"�W��;���%�[� q[����H3�W�.%��{s�\��@�*��˟�yg��r��#]���"�>����5{h;j�����8���"�QE��h��J,�f6��^�)|�X�]�bO�Ȋh��dZ`��D����e��7����f� 0��L��!�-m�r�md�g�읬��8K`�2(�T�U��Wl����C7���C���7@C&�5q�����j�gȼf3#�l��X!�/z����"�qi��{�8C����F��d�8J���pH�%� �AO�另�1����]�P��V'A��Țt�j�ba�9���0�&��[��4}Q?/��M�^�����b����+sb���ٖr�>PU@�	�xS���c��ٴ}�Sa6���]�̣���y�Yz���^��сWj+�r �|8z�C�yzf0�5(&v���]����Ew�)�H�^�݂�x�opK��e�� }Q�`�1d���eA�9#'o7�i!lr����7��Ǒk-���;&xOX"Z��~�����4O�A�2h".���wt�q��{�MRu^�	[<ڊ���!��(Y�n���C�dx�؆��&��nSڰ�%<�6v� �G�\j��g��/�~���(�����u
�0�/':a���m����i�-,6�en�@Ңm$�����X5o�"�緿���c��\�֠���ʨ�U$��}��-)}�@þ�݌�K��K�$�+I�̴��d+�#���}_��6D��$��녟l�}�JlGv���^����cMOɒ��?�U2��4�K[Q�j=H�K�Aaf��iZ�Z�m�o�7���	zr�G�?QRc��@~w����� 8��a�u����(>���G����Y�ga�O-qp�	8#��}ҽE��-̰OF~8�{�\P��x�b�"���Ce,���E;�1�,ŏ
L��"d1$(3!�ZB��]Fj(Gr��H�ߣ$Q��.��ߧ�1Ph#6I�Vb~�7�l��κ5-B�F�5R�d��uB4�#��B��������Q��؟���?`�km6�4�#6�F>t.�j8����v���%���z�/g���g��z/Ҁ�,��l����q�\Hs�����phmT ��-�$.[]Q�w����Z��4J?*�dW��&�x�JO���7��R�O Ck��ĖxFz��)2 �V��l�$9	������U���MO-ƞR��.I��Uǭ��p~i�*�wB{QsM�S�gf9R!,`_�9�Tq�b�w�"f�W��88K't���f����geg���Fj�9g&Z�2�z��3�N����D�n`Ā	�KF�AyK�"I��Cj#��졝�<D�Ź�C�Tt ۍ�oS����?��#��'آ��v!_��V��.��X"Σv_8�娟�K�CC
�zU��g�1gy��|=!h.��
�JZ(6����fk����ܦ�"��n��b��c��V^��`G����v=�3�}rI�I�QOt�t立|)GnV[��%��9
���rD���Zy��)u���A5S9�}��kYZ�22��럨��7N��B��8��1�� HpO�h󅫴����!O Hr�q!J�� ĕ�,�sJff�@YKL/%3(5,���'������
F�.G����q݄��o�si<=ܺ�h����צ��Mr��{Ɔ�Vg-]2�Ag���.v�1Ɵ���eב�^�'57H�����-��(�4)�\؂��Y�@}s��Q��ˉ�m���'�uZ�ʃ���T}Cs�ſk��{�~?�a�h�^���lp1H��E褞k�W=��5�5\pD>^�*�_�U�;f��"A��@)�{۲�&]�->�|�z�--�O{,n4����
Oc͵�C1R5�D8�W��5E�\!sǏ>��'���n@$/T2P���֊�e��}}E��O�b����&ȅ��%d"���@ �eH�iDVf�7u��+��n7��p�+�d3﷮�v)aέ�f��D��4ْ�y�ó�7�jP�r�@�OL�~�&fd�򓔎���x��ec
5�S��BV�~-ĪFm��_�P��MM?4	r��,v	=.��z�tٛ`"��6��D��ɰC�ޒ�Z�����ح޲�����;�����iM��D*c`��,\���E�֨����WG��B>�*��@̜
D�k,�m�������Md(���+a�l!�㗒�}�Ym 
����6=]�[?ͩ=--�ٕ���%y�FB|�氠�u]���1*ޣ��@���Dd���a��|�^q2�>�!�H��6��O(Ѥ���S�q���ά��,���ߡ�s���ۉ%���U%I�����������ƥ�s�z8k���+KJ��;�A?�V�������+�r9;ˍ�Ęx�k��~���Y��ȵsg��Bd�,u�DF�܏{����P�s�����e`����Ť"��\���?aT��<�U�V��B�}��+rQ�fkw���L`���<�iO�7l����������18�L�@f	�ks��R���#��a�Q�>�+am)J_�P���xĎ2τ�dX�;17�V�܀2u9���k�I�SC?��O�b܆��Վ��%;D�s�kΟn9Kj ,.8q���u_�;u��5�X�B��mP�7|���h��y9���a��c�w�G��Pj�_x5J����If<�H�:n���1��y�a|e�
�*�el�z� �e����OpDe��F�U�ᵩCJP=�����9�B�e��c��,��x��Y�s�-o�Z\��7�Ʀ���T2�=���x{8#�"�-5eΞ[<�ѱ�MwHC�u�X�hR��ޙ�p8�f�s=&\�bG����]��<c�٭�B �]W��lL]~�,�8����ܕ��������1���U�c�:�[�w���kл�`H�W�b���F��_=v %bpֆH��j�!�� BA�Z��of�e���VЪF o9":z!	 �קd~���b�0y�:��:��ܯ�҇oW2VxS�y��a������{Av�4��n�Y�A��Ix�d�l<N�Y���*�p�-G+��Kǚ����.�k��[�Em���AXfw��F7�`X�}�
+*��2;�근ТiD����I�QK�F�z^�PFX(=�>��f]?�!Ҁ���e>:v/YK��DR`��N=F�d��`�ԳSPy��Q��ii��)�)��d�j��WR5�S_��e��z��6��7jv�����@���]>G��tW�	�[tc�X&��� ����rfIJI��#pM�tk+�uG���dSp����>8ϯx 
D��==��ZՋ�vƞ�Ȥ�TB&0�=��,ܵR�������5^����dx1�<u�)����	l�f`o�o^!�o���e��^e���s��\� �Ϛ���>e�Ϛ��9n�h�f�/٘�[,���\[y�r���?��&�CN�����D�0P۞4�y�G�\sVH���-��m��&�`�}Μ9P
{8��C����&^�L�2��g��P0y��2�Ra��`�Շn�ܓ#�4{ೄ���|��!�q����'m�?�;[Z[�i(�ߍ;� !���'�m�H��nV��Hq!
�_{o����L]�R��n���>D<����:L�0o4+�����ҲȔ/��>Y�`�}�	x��.��׈UD��_�S��'@f�b������!���x����}Z/�h�iw��a�%O1u�5�e�>� ��!a941�lD������6�ڜX��L�X�o���6�$:"�Űq��5����z����Ɏ�A�k�s.9���%�N�wԸݞ�e:�����Yhy���$&4����9t����ʷ �fD���~_��Z-��1iA��>1L9��M꟠䬲dq�H����F���jy��g�Q*���(_�s�cJ0���)��i�B��6��z�:Í��	���\�9˂����˽7Q�:�!B�<���AK�F�'ke1�5��;���*�X�%7��dd� �Z�f�x� �����!T˝�]�>JNϊt�?q�ߏ�OCC����Q����߆LV�տ�V�sg�R�ż*��$3�ߩG�����?O�mNe*"���7D��{ś���,~f���IP���Rb�%�����i�M�"���.���S�1����l@t;H�Ol��Y�؇wh[���৴�ҁ�EK��i�6m;oPw�ʮ��큎��x���tk��N�F�!��b������Z?}����E��q��tѿ�J]�"㭈E�y$���û��W��O0Xu���T����BpLflc�6�?�^iF��g���PFp)¬�~�}9�啸�/t���qD�U��uI�o��|��5��;�,�3����Za���O=�a҆"I�����u����v���?��(r��R0���r���54Y\d���D��Έ�V �0��ƫ�]��T^�	;է���g��n>Fɳ}wc_8�҇�:V��^!��A�� �0)a��J���+��i,�С�d7̵/�<?g;ܥv�7�U�