��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C�D�}U(�}kz�����eU�y6e���>���s,�p]�$�$[Ke½9^E��E6���9�Plo�(�+����`V"��!�ma������x_��RF��|��\�x�p%�.�47�ͦE��X�;[�n3�[oF����[xZT�����w�S/ct�h =��~"<�5s��N9��	q�{���7��]H�H���Ċ ��?5�^P2�,P9uMY�7Tv����m����_q�>�}'�V  6���v#؟�7 �o`Iw��%:� ��jZi��2��O6A��`	��P1�Z\����:��ekBRwEq�ĥ��5�aQP�pw�I���vH��G��z���j䗰�Ѓ�M���6��u�N���X��+Q-���T��:z��W�ۿ@K���75pbi,bTފZ�s��րΠ�L�̘�"�F9^�j�p�oʜ���P��	���|��O��Oǂ����Rl�R`[,����@���t���ά���c�������i=���1�lffGl��.iP�/�����A7���O�|����8����Б+��H�pQ�o-b4���R�d<��*՝	��Z�5��N ��d-�aK�J/{dn=��9�fz��-�%U-/�D�D��m�����;�*��2%��fZ|��&��B�>d�{��W��6foJg����0�̌���������+���tfI�e��P����/'5��s6��~ 12¬{7��,�Z��~�{&�B�w��.�m���0������p���X����"	2ca�AO1x�j�s ch���3���'�麹F��R�;X$8/�`�� �Y�0r���览�{��]��}�T�l_ݩ�$Tz�$>0�,�y��XGb�