��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V�� ��9��[#��`�՝'�5�:I���A�YwF��PN#u��Ts@ϣ�/�F�`@X#���R���Z��m9�P��dxt�N9/�=��l���}�,x�PH�l��n���-��j�%�mĈ՗�[�^�Z��0%B��(^}"6QD��|h�:ǲ��I��MD�8�Z^�H�;x����ޭw�L+�.�G�'�!/��}fpB�A��m�M�A����v� ��;s:���A��lTN�l������t'��\J��ԙ��ϐ��#YOX��<�}2�d��`Fx�bƻ;��k��`�&쟮��k��F�C���8�69�l�%[��W$F���*�?�P�������7��AR>��!��m���.�c&�2�#�������(+��vH�J����pB���ܙ:8'��T����A>��}�tV/ �dQ�9w�ǹ���ArK|�?�U`	�����V�m��Ήa�M7���j~��"U`��N��1��`�v
ь���Z�c�<�����7It������%�w��QѺ���V�SjWm��V���r΀�mz�z���#K�~��_u�������TySJ�9a�	��(�E�X����e��_,��[����o��Rٕ���-_���-$_d�����w�d�`�* �Cܛ��E��k5��9B4���W�ä�`�-V�pǎy�V!v�Х�������J�E-�yV�&�H�2^S)���g����c)��X�������w3>b�Tȓ�P,�X�>�(Ϫo6�m�x.����E����t1*��J/
�y.�Dw�'�Sl��U��^]ǕK,���r��>jJV��&01�D�b�9�G´�zҮ���ܚd1=,���p )�g� �	��9��o����������{f��XJRY��eI"���O?��+��e�-�'��MU�;W�Sv�b��j�Oi��S��
xp���9�����5_S��w$ƧrdZ���P<�:����~H�Rt*Gz*c׽9��&I��q���阈P@\�����m_o�I��ĿRh�$q�I�o�[����Rb��e��:{�Ll�ZL�H� �]fh����dOF)���m��W� �b�Q�߄kqO�>��|˵I��9?q�v�j�u�^A�">�~��.u�3{��|�5��'r$�M]����`i\�{�����*v3�X|Vl�|N-XT��@������!�����X�^ʹz'θM
4|&%��+����FE �tË��#��0(�MH�]���ȓ��d��A�i×j�3���@�&����>� �(è��τ5�.�Mw}���U\Ǥ�m�T7*
:�WH����su�W_Tܶ9��h���ش�c�3�?t/���r(���"MP±^܃$sF����C�}Gi���2��.|����A��ў^����@���6�@W��5��wg�L�4��#���3T;�Opk4��2!����̵�_ƹ\#�B�z���D5w�C���K��AC=wЄj'y	j	5ύ:VS�UM�g����e����R����1��5G�X}���L��)F3�`E��FeV��0�G��e�q�c����C��&ː��/Z���ʥ�����Z�8�Ql���q���}�,�:��U���?H)*����o�ǻ�v��0�T$CZ�� �R`ۥ����g}O�^J���Y�՘�_��y;��3V�����\��g��6Gt@1�]��l+ =��y:�@�j)�D����D�d��Qao�Y1d!u8Z�Ӭ�aץ�U�d�t$� FH�5qJxWZ����"�E����N;e����Jn��|�1-�7ˊP��ʇ�k��,Jվm��+Ku_���0�a�U��H��w��B>	�E��E�aE	�VOa��D�D�[KxPZ}D��3^������+�f�7��Tq�Eg���8+�(D��R�eΝ����ؐ&�� �'��d�a-�HB��d[��3�;i���P��5�P|��
�4/�Ը��#��@��hJy����E:���j����o��ѣ͇�H��pqv������p��"k�a΀E]˹2l����s�H�h�VA
��ږ4_;0Vbe�u坢oV���w;��/D��ב�N�s��PDShS:��H�/^s�]x ��o��ȴD�&�u��(}�^͉��n9�mD3\Anzc�����K
$D��48�U��e����;���A|.9-��WP���'	��K+�ˮ���-��i�� ��UM�Ë�j����L������\��U_]�q
^E����A�O����N2�	�~�ʿ.�<�%�'6�����dͰ�x�	�ݶu��=�����)��J��������2MyJ��G���{V.̕�����ǘ׈c��<S���r� T��6�gs�\K�_V-m4��M�}�}�ـ��S(�n�<\d�<�wՅ� �sT�k���"f8*��8�K���Ņ��$ϐr ���cp�g�����g�eg�0�iIkt��L?{�kbG�,6� ��Ǚn��_R���Ec�O�!Y�zvAB2Wi�ҧ� �,.��.�W	t�[*�9X��kx�JX}g;�7�di�Տ�HS���a�D��;(e��}�y�4q4B�t3B����0$	C]�'�y���.q1;gm}�">�r:�I:��o-"}�H�A!)��4��s���%�O��u;��~