��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V����hN=��a���)�硹<H��׮��`̼��D�g�;�mR�#rj��S��k@'�q�/�ha��pc�R�(��g�F�ו�����`d%D��G�qK�DW�+X���iv�O�O����9�t�0���`�<�F�2MGJ�g_Ю3����Na/��4-^}��ru1������>�9��& c�dN���(�lE#�)�<���4�z���V���i"�h�7�������(J?�⿱���~�t�y�k�)V� 2%��ޡ�)Di�6�Xt ��p#���D�%wS��.����p �.�U�e:�ȓ#�31Q�5��q0dp}x76j:����MA���0μb��TU�	�iwNv�����ϟ�J����T?�>�8c� �w��@�( Rh��Ӄ]慱ݎ������*��PY���[bp�g�Læ�Es ݏ^��P�v1м;��f����$��s�jH_~W��:׾�>��KU�%m�c��C��e���x&�[ �g���JE��2�� �
"�k��"������~g~Fh78��Zj��7�+��E�8���Q0�ןՔoę$�D�,�s�,�m�v����x�v��2��{�E�VN��i>�E�f�'�6�)����h%�s7q�s����yh���i˦
��Q`�M�s���&���[��`I����g;%\�H]ד��ku
�(�����?�.E-<��7�o�!�ϡ��pQ @)�	\���Iy����>K�*(�s���I%k�]�#�����W�]M����(�>e� z�S�d���yp���v9�(�Hkf�'��ɪF��Sd��53'�I��F����	���+�g����5	�7�-+gdA��'�Aǹ�o�.6�^�˴��>�R��tꜟ3�:�r;��<����.��⯴��H�ҩ�8�x�[M9ִ�	��Ui��Z3g�	#���"1.k��;=07!�֢>�a�O�OQ��}�А2%#�Y���^>��"1qw���ڈ|,�|⧔ L�g`Ɣ�%��~6o�M.� ӯ-o%�͍M�<��*�B�m8^�vcWO&l�B1�,�/kT�Ĩ�h�i�`q� ���8fW:̞r�/�î���E�b=U#�H>�<7�'�)�!bC�y�q�r
yՀ0�I�Q[�zf����n�gL��b�I\���=t�@erܴ����G�>�Ýy�4��J �(=~%�m�T{o=���3tMoHn�x�QJM^
��>؍r�w	S���ܸ�}2��Ԩ�?u��t��رEU�X�yK5�E@����r����FT[ÎD�\E��{�.��F�v�<O����G��h�m�'v5Hn:g��x"7�Y�� "����ٴ^�~cǏ���ȋ$EF�~�YyT��H�J���߇gTb'��ZO�E��֊�X�+䗿����ȫAq&uB�V5�
����ٙi�֙�Xn#A�Pى㼾L����$�
�垠��7|��	H@���7ʱ���3�
�N���M�19���=���ek�OD������S�������I���io�V�r.ь�<B��Vd�C�`�\D�c-�CpO@�5�y$!l��V8�@������c�s��B\T�����n�{��c��pwM�����Ϊ�d�����X;D/�ѩ�ս��6�X�yn���鐗g����z�+�����|�����,�dJ��bLl n9�3ӔX������JX�S��s+���/g�������~��)�r�X6��q�'7��'^��d�	N�jH��ڇ�Ѡ��09m�`ӻ^��U�ǟen���7}��#��֔O�^�z��6�E��=C�T������U/+G��&����2ti��Т���%Qޫ�!Q�.c��a[�lh��Aَ��'�^�L�����k�a���#pQr��C�u�͓��r �b]P5�qQ8<��{!�Su?0�ϙT}a��K	\��WE��;���pz'��v��t%V�A�X�4{�KRG���V�s�j�R|���]�?��u�]��ak<���IK�e�!L�?�W{�o҈��;]����S=���@w�b51(�+)n�HW��!����q��D�S���8��1�i�jdV����Cxs^K�/Q�Q�f&K�P��_%�*Bm�M��o�V�7�0<�Lv����N�_b.r�s�>f/k�K�[��ܮ�r2LU4y��%���?�t���^^�Y`���mRm�� c�Q�Vˠ8�YXB�f�F|�W4��Ⱥ�Lf����c#�����B.�9Sp��2#l��\��>ƈNCg|a�Z�M�7nO��Ė��\�R�F�8�gs�Wp��]�z� ;
�����?\<7�ίġ�K�!g
4N��!Z%4�*��9>��L�����k{��`FŅ%�m�Q�*���rݏ��-�^-���B��N&�!���B�;�m `�1]A���o &$"���{y7���7"g����Ւ��kS��GO&v��d�X	/�r�ǿ�j�S��;k9��*;[4��ug&�2�ڽ%�e��b�����!�l�V�̍��,��~�ڳ?8�]Q<�r��۫RW6�]����Ȩ	q@���:�j͚���5"^��]L��R!v{ �~qƏtv��Ҡ�3���&�4=�z�6�6�/�U�3�ˎ0)H�L���"D��^{�8"rR �H!�i���ߖ�f��`���	��XZ �}#S�M&@�k��f!��ɻ�߆'K^g�g����5��zͺZ�y���������<�8"o@	��=X!gd�ek�tX��U9�7�>������_2�A4RT��eK�V�Һ��=�Ns����ΩC�B�	�|���ۍ�o�Uwt�7�� |s�{�#�_jc����NK�32Q��y�Lr)7�6`�5�C�!���&?r�j��WCce~�G��w��=�م�Fpg����(�b���y�煍����x�+�2��Ɇ�ұwBȠq	��=�iH�悗��y�z�T�`�/���kM�>���	Ssp�3�h�p�#T��	n'���6�+9#�y���ue.�A+f""�4��
L�t�M��F_\���v�ҽ�$���������SB8q�<L�7]�����1G��i��&�	�g��(ӂ�"-V�:6y� �QMB(�#�%��N�`U��)����}����X�|�d�N��}��cX��(f^���/�b��Ѻ��XT��j
��X��_����>�������]˰E>6?���]�Z����8PHש����H�u��j+�=�&��8��GO�w0�]s�[��.��Q"8��z8�=�ѭ���fΰ`k�f��<���?[VtK忽^3(�ioRYH�Yt*,+Ut��\�o��J�����X�h}Ȣq�N��yt���%��{Y�F1��/B8�����k�Vv�Jo�
v�=S��(� �o��t����t�Fc���1c�Bznd^`�G.b���ZÏ����;�n��|7�֦���x�;N v��A��-�M �m=	��ַ��O@�Z��Β���^���R�Y )��� W|7&K�f���%��kCЄj�sP_�k�זּ�&Ҧ�OS�t4�V�=��!����Yzv�m��ZBdllQ�of����#�>�ـ�Q�����϶�t:L"�ۻI{�8ےg���
��(��n��^Ӣ������k�8��V����u�3]��P���̪&�d�GiK+e���mv Ol��.��W���<j��L������ܸ ��{m���<tG�X�	���&�|���w�<-B��D7֑|	>F�Pn��(�w̌���4�C��'�M�U߮����p�#��rkҙך���n�Gg�ZW-���Y���d\�J�?�j�[aü���- >Eā�Z��Ke�s�<�޿v�����K �Þ_4��}&�֬���[����O�Խ��꠯����?���q����oN�# ��<����)�8���s�N�X(1e�6/���|to{�3
��Z���Z�Q<=1���^���v]�yk��vq����%P���@T}��It��?�!�k�]������x%�BRtj��"ۉ?�������\%$ca,e����?��ib��̱P-�`��+��\��*`�"ţ�[~��Nވwl6=]Kyp�G��q%�Ċm"��8ld�XI"��������+�?���i�bxeU�1ͭ�pU�����
����d_�$:q$�r�s��Ϫ�������ʦ>�L�n<"E0K�Ƅu�jZ�{���\���*��<�o�d���<���Ƚ� {؛��_SQ�����@I�B3�'!ۮ�0U������i�ї�}�j�W�R�������AUs�w<�Ck]�����ẘ4?w����������t>�;���;;"�ϔ��s�m�m�y �lv�m�%���U��m����S�L�x�XX�V�j+�{��@7��iYE9Z� �������H���+)~TV��@?9��A�g�>	���	��^.촒ڕI-4�n�Sa��Y�l�«��J��JJ�im�	D���^˔��*pjx����T�gލwJ#|���q��D ���a�v�����T���E5�����S�q� �}r�Sz&3%��-ɂ��l4��5e�6�T)S Us��X��1x�@g��s���*F�E���n�*�����S!����?A2��g���g�?��@'q�Kq��[�)��q���8�C�^���L]��"(A§��k<$�Xa���a[�\=mm�(��Z�X|=�!&������y:6w+�q>�v�ѻ� ����� ��`[C����
�x��:fe4��g��5��y�9�Frw9��*�Ԃ��s��4;�G��~�1�l�� Q��q�k�ʊ`EA4�r�<"Ǝ���>�R�B��}W�XEBB�}{9�tM�Nd(pD�V���+>;:*7DI��l��[b�$\���0jR�����c�����B��s.�"�q���Ũȳ8��D��C	�eY���V4OK@TЭ��L�2������ن!���b�XnxE�A���(��o^����j!"'�=��.Z�@���%��"�ǐM��h�Q���_�ʝX?��r���I�[5��t�^MáMT�ӌ�Ù�8����yH$�g~�v�M������b���^N����s�DZG��E/λp�^fQ��O��I�ߧA�}j�%;i���������E���5�0���AòR_ѓH��A������?'���?���_��cȓ͹fsM��o�8ьQxB�i�ɺ&�^��j�y�D\5=X��j��-���oV�5��h�Q��j.�-���l�SOVj^Ac;�uf;-���*��E��
��a����>��0��u�����v;v�+����^ ���0Z�����FjJ�1�oWH��u���H�n`�m9�뷇3Zj�ȹ�5#x���u���z�`�6:g�'tP.Njo�{����0�,��J`/2E���4�n�)�d�߄������S�o���#u��� X�E�5�`��s���OaZ�:�T��,�"vO'�b6W�e����(������l���EWJݒ�}K�?%x�1�:�,�|�PT�q�ʊ���~�����K���c��p�/Z������Ob��Z�S�]�K���]�	v�^�	�f1�5<���aΏ�M^��S��yO6��&�������k� "r&�f# �O�rԌeg�M����}��3#�#�d�T��^�M �5^��D�nl�]�\�#<�O^��>�r�"�l
'�3'iz	���Q4\����p%o��G����<�۫"s(c���m�&�K�-�&��o�a.L�a]���PӬ�~+p��e��&qvSJ>jaj7�v���Χj�m�h�:EN�mi��\'���3:�ܪ}
�8dz��\ք���1I1�A:�=��5k9�ں�0A빠
��M�_���6���P3�mޗ~<]�y�|l�k�P���C;w�OAa��}���)�r�f�y��2��?��>�k���d�������kO�ҳ[j���)�^Rʵ���&D֑��a�: �m��Lyߦ�w�P3�2U�*`/ڽ�廹@煀*�%�R�Yt Y�M����-!�S+�v�3�Y>�bU
�@@
	2JD�>���-��+⋜O�]I�U7e�)��i5m4( �h<�%�g���|��+�(��<o�*/����B����=�c$���xeE�@nA��MΙ�H��YUOU�R�{F���V�o}�ao��	|�4X�	��ly�!Zb�G����(Wg����6al~�i�=��Pj�I�ɤ5�����p��x�uB#V<��:��������v�u�W��5�l��ff1�f����bv�H^�*�����Db^Ӓ�xc���7���5��V��d=3��Pϯ�d�@#ʧNB��(�.�B�lا!�wm���?���wP���˯b.ˁ�����8�/g��m~و��8�m��ٰ������30,�<�p�d�
v�[������	�Uz!k�!["'���6]�dcҲs.cvO'��i�>�ڜ�ګ�+Ģ?"	Uav�)g�L���h�Srn�HE��
��_DQْ�W$v��۶�)�ɜ� 0�'^��i���O�ʵE�P�LlF�����|F��*�U���@�*Cm�Z�"S��eν;�fnk-���6嶿].��;>� �󞟵kP$�x*�q0�1�F
��繬����DV��[!��h৸�&�)Y��\�f��Z3���i�T�ȓ��h~��c1�ݍ��4դ7�h(��k��sV��i戎Ib�8�%F�ZcDQ�԰g;X+����l9�ݫջK)A>���B��Ҡ*���?��6�Y�e�|Y�S�)�����F�/����g`�����la�*N7�[�� ����c����<��D�4G��{W���>\M �sE��Lؠ�3P�w��)�ϵ;5{Z
W���6��)�n�M��v����Y>q|,n��]J%�U%\a���6u+0Z(�1,fN��-v���D�lA݅4>�_f�O����2��Z\��Z,���B������r,k}��� Yș_�R<��Pjy9E�X������$���q��Y_�K�Mh�G�B^`�#=���[�ha��Qܧ����:�����ZOi��{����wA^��oD�4|d!B(�J��>��o������$7�JO��t����s�c#|��("�蝞�Z�C�,:SA>8Cʏ4T����Ä���+ڻ#���l p���\e����5uP��������╷�=	3w��#8=�T�U�k��^�=F�eB�ew���n�e�WK����T}�OD���M�O�D׮G�鐸3Z��v��� 7��
��m��&b�����=<����LV|�w����q�����A�^��@St��򘦕9l��U�3�Z�+�Z�3��Kv��4��UY�&�ﺇ�U?)�����Tu#��o�S�:q?V�r�j���13� �p.��X��N��>[h�p���Qo\ɃS�#�e�#g�n������Ш+�@��А�V�Z�Tb���BI��W���9�5H��j_��l�g~"��@�ۖ٘�Y�4ݑ<Y���:$l�lT8ԭ;��(Ű��g$���\e����3� ��<<:KƝ�d�����319�_���<U�@�-�4f񈗼a^��*�M�Q�W=�����(��C&��J.�����SQ���4�"��i���?����,�p%[���7�������qW�g�Q�:�t�.Tb���X��;��J�OA��bS�c�k�gG�h1�,L�9��D1�a/��s��&yJ�I��bB]�@���5��e�j�� �傗_�t����~H��	B��m<���U�ZKf�Ԅ�pfz{���J��5�$Eo�9Q�Yg�T`M���2M�)xR�kg2�Tq`�ɖQ��k,���q�t�2y9�my�ȳ���j@��فB����/weoq�	{x�����c�fZ)/ A�9����bk{��,|�	���}�"^�۲*�o�R�]�r���T�{{��� {0"�l@����/i����DK!o��_���!tY�j9���7�b`'�~o %b"z%!Vl�Խ��*s�])1z�v�Yg��$��<�c2�S�@�Ѱ��y���;u:�FA�htb.��FP3�	�80N ��jn�)ÛP�e:���җ�v�E6M�)ڈ�m��J�������R�8�iZ�"+��Me�n�[[�-I�]�2�ݔ��,Q��>&&ϵ��v�Ʒ��N�C|�=��
����"B֔�'� 3��n�	dv��B&&tbY��X���P��C3�c/��\P�g�ؽ0	SvD�B��o�dٿ�Q�xy���o��|x���%&Z��YH@&.Z�=9��_����vǻ��$i���o?��,��D��y��ź/Զ���7z?��e�����b��?'p㘮1#���@`��c̓�>x���V!>��DX� "9B��O�t�.�FL��[�}`�ԖU?�,@�Q#W1��U�甾U��McBU|S�曂�Qxd1�(p���jm��*�^�7�ʔ��J��SZ��{5E�'"��D�Ʀ�-,�^}��_V>J��ሤq������F�:p;l�����޾~�O[�)8�i�it�Z`�kZ,�7O���i����n~���GgL��}�f����`�G�)�#���[�s넌�V#�?J֒3��c:��զ��@��,��4 �Z�	���������[6Xtc��j�C��2&3a+JNG��\����r׳D�3*?����j�x��5���l��Վ���ŭ1I!C��r٬���H�TF<����6ߩ��l=�L�kׇ��W���E�%ġV��b`*���I�t�,	�V�K<�B��K�a�N�Z`�Z~��m�n,�E�v���?'u-�'�a�1��.qp�6�g�g���t���/D>q������UkO��`eػ>l��^��B��ʪS���9��|��S{JOu���(��0���C���rwB�>4�+?oE��{抯�'zi�i65�
=���;�A��J�[��<�o����U7��R�J��*���#MB(:h4�E_J��ڄ��;bxC"~eF溝)ҏ��`l�t綞3��J(�Zp�A+.�Էyf�#��^����lH"f�t[�Dl��2[Dwl��_G�MQ��9i�����lh�|��w��c�7)5t�s}�P���T���3Id���ل߶����-�!��i�a$�ܒnN%-�Z'��q����7�IS�"lV��IɩΓ�t�Q_:���'#���L9W������������6�$�<ـ��nsD䃃2�KBZ-�����S�w
nQЍT�(����� A�M_�4�h��3�C�qv��A U����
Erϐ*J�loTE���sRߍ顱�)<�h'؋{��z��H�'&d]k<ᢙ���"v\����PZ���bC��8ۗ���ǿ�l��П�N��z��S�M��&t�X��Ch�
Տ6�@�+��e{"�7q�#�K�S��R/���OV5�������,ɀ��g@���r�B#�x�w�&��F��д�f�h�Yb��\XS�bV2R���0_�Rx���s7�F�����L?��u��/Z�u�I� ~�~��pf��]g�T������p���ӹ���910<^{�+����P_`��aϬU���0;�+7�Qp5�}N��ӓ�����mvA�O$����������;����ۧ����/���k�VP�\x`gPE�q�K�\�I|���?cl@�5�2̻By�s��k6L��=ogv�p�x��${�r�+�_�D��C���D�e���aB~d��3�U�o4���3�3��		��w���z���W� ��)Vyj;�sI���Q�7Xj�zv~%��X��]9���맾�.�����f�S�;�'���.U���Ѩ�<�bG��>~���G��l�4lqbu,L,�|��#CǺ�F�ѭ���p0��s=���"��TO� ���N^`�j�״���Pw�b@B��W�ӂ�J��-�����(�#�u<�:&'���f�FH}{*2���7%��������=�9P�KB���t���A�oD��Y�4��?w�ԥ���W\l����c	�͋� '���������^�.�]�R�/љk@��@�7���Id���Φ̪5.G���D�qP	�M���T�(�h��h��־a3�pIcu����w�P��Q,�I��wq=]㉍���CG����$9)�bL����?��zZX$T��Κht��A)N���榷d\G��`���79���:���I�C*�6�BIgC֘�,�n�)��I[�"Z�n�o�2����!D�����"�é�� �G`�m�T&�Ǔ ��\�`Q�6ˉ����\��0�����(�%X�ԓ�.�ٯ	P���؝jQ�7�-�Uׄ�IS�$P0K�+��>��̥�4�|DT
n���TG��(D���&�*.(�=y'��ʒ���!�Z�Di���YW�S���ν�j��(���`_��&�L�"~��?Tb���,Lc��;&%M����R��������B���r˧9�/�Wrٵh���~|�a�?Р�������d��v)�j�w�"y�?�yL��?�r
�|B'����ɂ�B~�!}��ò�U^�aq�UB0`�-Q���j�������~ԓ���k&4�׏L��c5���ؿF��[D�|k�_$��Q����<��	��EP$���W�����W�7�"��A�"nT��&M�xLC@f5�[�Mh���6�2S$����9h�lJ������c��������{��\D���Y12u>d	V�cl���Z㶒�R�T��װ�[=j� IFqEZ��μ.��Jf6�{h��2z��#��*�h�Rt�l̝��EK�)F�}b섆[}ƙ��A��]ar�#��&���Εl@M�]~8��f�D�����?�C��d5�]��r�[0�iw���cLF���)ʿ󓩿Ap@���N�VF�I��~�{�)�q�8�!hw���}Jr~�}����!bV��� �3��F!�|O�`bw&��E�Aw�B7��>q���M��GV�%8.Y�n��6��h+��00�?y�g��c	0Ɵ�%��0�j=��إ+����j)��_"o|	�V�ml⨢a�R����Ͻ�áYJ/7?p���6�.4"$J��<̈2p�5���D)���;:���)Y��D�Jjc���X_��
�wqXCZ��b�Nr�9qc�� ��a�ݶ��2�M����{��/�m��Eu5h`���1�p�;"����kt��Ū-�Y��t!P��&N �?p�Z�X�@	�����_N5��P�a���s�!Y=)ܛ~�+=3�0$-��)-�0�ᥒ����hI/����AZ�����������ۧ_�;�L�^	1�B���D��EV�#���n8%�}f��+\c`��@���ȑk�㽫�� �������CgX�y������Q��GZ 7M:� �i��3�ٷ�{o==x �)��}TQ� � e�H�~��.������ϩb��,�I/W�P��lF~�)�[ۨf�Y�/�z��>c��?�й��h��8�$yB�[*/�ZEI݋��#Qʔ�rR�诧nB%�5�e$x���`�
�N0e�a�|V�yt�]���tAkQ��f�k���;���P���ს�d۫i쓯n��5�� 3@���A�=ɝ�1/@<��}��"�'-�t-�JCH�\���a0N����]IM��,`{��Ĉ��#A�xe�Du���e�-aWmU����J��6,*F��p�|�8���&x�ce�u�[s[Â���ս�����f�(2����Yݨ�o�0�����+8����@�V���+@�jVs�g��'���Hnb0<�hs�QI�$�8�[�M0��2��Y��P"�yCR���Ge�W>����j�tLC�������xHQ`��Y����ũ=�Gk����}/_��?���vJ��� �B��0Ll+�t.�h�"ОB��X@Rz�H1_���ki�(���}S,�~ʼ2u� 9���%�� �L�x����o'���-f��NFy��T��<nG{�O���madMU.Tq��Y��[��V6�z��1�&��R��a
'n���k'֖H��Q�m�6��'�k���.�o��f!F2���7�d�����>!e �Q�ꝉ��6%☨�'`_�0���E��F�k�M��Rq4�a;��=*ݖ֤M�!]^@����+T�԰+�a�f=�+���m��)9`^�*&4��4��?�,��[���P�"��-I��*��e( nQ�8�1���f����2���%;P�����:�����Ƶ�e��i�)��_3�A�����]X�>�A�dWvU����5�Q�Rxib�^E��{��)Lu�7�Ak41�(Nb���g���|z��WV��V�7*�鼘�@z�QN�I>ي�:i޸�fpd2�)�|�C�9$�M{
�9��ݹ�_�����&��d��z��9&���PP�d�S:O�7��E�e����gjY����	}���@0��J�+��:=�m�#��v}����!�S�_H�d4Opf�X��[���U4�w����W$>�x̚��Zd{�_ްSS������� b$��㮬��0�4X3-�H_��"�djBv���z=��{,�n��]����k1y��(R=V�]�N���'�O|m^{�,� �&Z{��6���XrJZTy��q=�8�(�}��Kl��>�?G;ycRK
`}�ƴ�8�1�;D8���僪�o/}JU/�+V�_��!$/�,)�{͊)�pPfc�ox����|��31�s�7
f�AR0��K�5٧<T�}���:���6�D�g��a��p�Ds5���d��)�~��5֨H�|,���ݩpC�r��w#��q&�(D'*�~l*y���l�j�E"��G=�3f�tys�-�R1�� 8/H3��p�)<p9/$!v������ �\�����?Z��[�ǻQF� ���%	�j3>\/�n�=�c�۳��ړ5�%}�����[L`(�4bɥ�ާ%&���}��+��Ġuqr\!
-����f�o#��Z�]�ȃ�Eex{Vh����(iS���H�c���QQ#Y,ee��Y7Ys�t�0r��2D�Wt�c6
��u)�
ъZ�S��Cc���]-q�M؂V䰭�����(7`��S�qU{�����/<FK���ou{r�]�_D�_���|��#��\q�c�Y4J���vĤ��6B�(��}K�Gzw�Yn��M��U�ؼ8���t�|�`���7�x�yDzc�K���5}�7
7�&����#��

��;�v�;v�R��ιT�*�f2����E䤂͗|X�Gx���/"i��Q�(n���"�iSh�WJ\B��p�R��O-��3����n�]��Cq���:?\qʕ�A(s��_���8Y���R&� $���W�0p�ZV�F�� ��;9B*�]��Gc�R�ť��r�q&�<������$�źs���z��$�=%A4	Rπ�l�o,���r��ʗ��A����بt�/O6+=�O�2$FY�*'0���Z�ٍ���3l��FWhA��&����h��L�N<�!g5�8��J]+�f��@��B�^��Cj���$,w'r�j����wX��)�7_�`���ʣ??�f7\v���zߵUG�
�����V9���C��"���o���}S8ߠwg��H[��Ce�/���p���'���k����s�oI�Q�s<x��EeL d�iy�?�X����G8�llC󓉙�&G�]d�ZFV�D�<.��0�Yh�	�!� ,��Ʃ�ǫ�?�Q����;6���w�>˿ ��8#��[��ᤛ6mGZX�U1�[ڔ��U��	lDA��K�w�z�OܸߤA!_��>h� ��t���]������x��V��3q�]7��.S�!�0߇��h��?�ƒ��JI8��M{� u�Z��0|9"Vn ��o;���O0�� ��7�ү��m����FL�a�*ug�+�F���=�cQi����QⅮ�����o�7!L�(�Q��@�쳧V�c�L��O��-��˾��:�v�_�x�?�{�� �H��²�$E�Q'����9�N�V���]6����=%�W�q����Īj�������<@�2��+�rN)�l{�:�!��`0�j$6�?&�=�ۖ�3��.ҷ�����(����TZԘd�"^v���l�+l*!�GK�JgU��	ĳs��h�r��H^L�0x��j�0��Y�AUyl ��7��Xa����"�8���y��Y@�$M_�"�����[T\Wj@�nA9��j��4���[_]!p��@�����	C��'�pqTZ�.	弸�r���ٔ]�yKhA��k39
&`Q�`˳�[��Fa�9��,���-�Q�2S���o�&�a��iN�vkE�[��|,e?�Q�"�	u�|�7�Ғ�R��k8y�i��` {��u���M+hM�Ƞ?����i���N��d�c�Wr�Tm�lll�0�p�xe��y����&7����g�n������V�	��)�S�X����K�3�r�Q~�6X��&����S�)hOE��!�7%���h�;l_�R�T@�N�ɑ7��� ����bĤm�9���.��0��m�8��O/0Z�c+����d�{L��:;�,��1*X3�4�7�]�K�}Dq���]�(����?�IU��P��F�
��2љQ��v$h͵�)���c}�Q����9!�LOr��%Q�T��$�7zٱ�Èhaw�hI����_P�9g�N��*&3�6����
�2�_8*��6@��u�Pl�M.�� �W!�=�;❌����������??��J��J���N���5Τ�Q ���`�H�k�)�����HwwH�&`���vƍ�$V~ß{�d{"5b�_�!캘 {���3c^���HW
L�f1�81�i�ո}r3)-�/%ش�_���&:MQ�λ7� ������v�l.�I^��y�������z�8C~cU���t������u
f�q�2���i�MC�K�e#d�q�X���Ld*ӑ*�X��N�U���o6GIp!�w�@���A	ʱ�~�X����'߽�~U���BT��������^��\u�f�ûL�����0�m�z,�gP�{�o�7T�!Y@�`(yւ�]lZ�V�z4���Jt�Z��KÆ�JܶH:��~�֥� ����S�+gc6E���lڐ�|];*��Q�j���+�u���Ϛ� ��4R��r��)�G}K;�ļ[�J$G��s�r��lo}��ߗy�_�4��t�R�}3��b�-D�x� ���{ƿ�+�}W�^��2E�۩8��xb����7I.�蓳ZC��,�ӎ�g�d� ����V$9���`�X�����r�Oܘѹ/�a��K��K#���e�ȟ���g\_%�
�� ���}�0�7�y�UE-$����h��
�6h����0;�f���eXr�K���Km1���_=R�j�3�P�&�<�D������R-��������װr,?�ԙ|g��Im�,���ME[����������ڙN�©~ؾt����>v�๸|0�&�X� �}F�oS����`�Eb ��QH�m� H���7=�>��Q�H�����J��@�r砃�!O���Q�,��.��� U��=gM��5C��Rܭ0�}��*}r�~�C��F�Ja�B/��Jd!z�\��Ε�|��w�����i\����ȟ �L@��a�T��"T��8E@w����:�YC�}p�]��:�z�kb�p4�sO��8f'�o�\��ֲ�6U���0��^���X	Y�>�
y[���v�o��a�$���\ꙋh"��	�:JJ���$�C%Z��=�������K�7�Z��(�
IMr_w��{\B��#���O�$6$Z�<3f�rR*�;-�c�o��Ic2����3iZa��K,�5׍��7U��%ӱ,o�j��̀��2.?6S����+E�2�s���7�[g��VG���aK#��G4&H򬉈�[��p@�
�Sf���DJ�A�ٿ�X�CCDemn�fJ۞�Z����B�6�y�����K�ì�/�J�:/��_|!�ɘ�FWD*�����9��O�-`�^��610�v�+}��B��%{](�R�z���D�=S�����e'h�n��0}GZ5Z�O�����ŲWv�o�]���k�b��F���3sVs�>�Q�I�^�.9��mWH�p\�2z�s�G���dN1x�񢬽2�`��T� XZ�E���A�LB�tZ�|V;G�P���h`C�����ײ�-'u��}Sk����h$ZuN��I�����\��#(�� �;#�r�*�\dF�\��Iv3��ʩ�W ʢ�/�3LD^1�T�[�۲1Yz���Q��=�z7�o��Yd���:J�kz������̓���gvt^��+�;XN<>�� ��dn?��_j���K�[�S/�70=�ii�Lr�H�2�C�&�&2Z�>Z�!��Յ�p�����t3���*�3��c�5F��Ձ+�v��Fp�c#�I`|_��!<�:��-�����9�G���~�+$�Hð�KG�$�D�� ޕ�;]���QֵN�V��L��ӎkX<l��z��Y|5�Z!����!���}6�AgP��w8�������b6��%�6lP�p��`�)���	��-z뇪Z�>�@�=m��ub�D@���g����w���g$��Q�K���7���S��+��+�!E��x>�>����/���eS�-�ʘ����k[��$IJmo�X�������f$*�����Pj )d�ܶ���Ł��Ką Y(�*gG��}R!�B�#���^/Z�8�����2J�o���Q�����o�n+C�иH`��,��T��%o��y�M$G��*��G���clȓ��mI��zKf�G�0�M���9��>�S����G((�\�;'g4�0aO����Tǎ���k�*��J�	�"�C.ѿ ���2��w8�b�'G�q#�e�|Yy#��,O�p�<�|̄T���9�1_���&����R *�$��/����T�$-+h�-����ݲ��(��j�q*��
���۴��u�T;6N)#�~2�U��&Oq������!5����8+�|��2	���k�rl�X��dak�,p��x��o_��8�D滱]˘T%oz7����0���iϚ̐Ռ�� ��Րc8|��N��@ň���At�$��tO/��]�����k�:r��/<���JL�D�����d
Z�>Y��!e�FL� �Ԉ�(��R�a�T
%8l %xZ*�����Hx' � |�B�nO�����Bj�;p��ҦO�M����z�a��4n�x��/j���7�A�>�g�X�2Ԛ��]_1y����+<p˧\-��Ei!��[..�:{%@1�3���v����+K��:Ǆ�:�pG$f��*�SJ
��NML�V�(�Q�jߠ�)���Y����K'�S)$~覇�����"�-��y��1�y���-����j
ӱy�Oe�_}+>v�?�E�(Yt��a��"�X���c&z/�̨L��r�I]�X� �h|'�I�7�/B�NQl�PJ$;���〩�������0�yG4gG���J'�t_1�Ґ�'Z��ƙqn����� ��$�����ʾ?3�e��<v�CS��ZA!%4n�؅�E4(e}שT�Q��)�� "����e���f�K��F��;+th�m����Gc5#�z�yH��]����?QV0�2�ƏB�L��N{�,�����n�!��3	i1{a|���'�����k�DdC�^��U�^#�fW�b{�#�+1*��]�E�W��qA�����e
6%U�n�A��W(ҍ�`�佩��o�F�US�<�%�����v�H�l��lh�$���B ��u�iq.��0�$XJe>(W������PSv-��G��geo���p4��Z[H��ϭ8���`]�q�� N��{���N��)�f�.F��+BY�/���W6b��w��>fBs�h�j�~�?!;R�)s�9��s�ZV�A�v95r?+.X`��u�Pr�e�R*�uQ�x��y��F��0����L+Z�S�uz	$�!�޷�(N0��W�A���V�x��1�I9�K�\]@ޏ�QD����0t�ԂC���fH���X�eѿ�+�
_���q���O�v���Q�g�I�֊N�u�~��X����r1�߲�=�1H8�M���0�\�o?Q��;�@�w/sM��
���'�sB�o��Z}�û8pq��8�	M(��~�L
�qu*`h���0nȨ�jM4�BS�rő���]'��u����]�(�[��8�_n�Q�n��W��xQ���ݶ]�jj��lL��?�9D %�>�@������ӄ�w�d�>���@�X��>�GE���C�<<;J>�D��R��74��&�m��
+���L"O|�Uf�f�lݝ�{����
���n;^���uX�w�¸LU�Z{�d���Ҿ0噰Nb� 
�`�akX���x���ݛ~G� �B����h�#���t��7���#����}R��Nݺޞ��ƚZ���{��0�:!�7ptf�M�aY���q�z���tc�C�CT�WO��>M�K��$�0��)A���t���pBTL��O�'.R+���[�W�m[4����8�i(�N$�Ȭ#C�޺nOƲ����cF'6(�V3�������3_��WW?��U�K�,���7~ ��6kH$�9�p���s<2354�g�e�E��֕��;��~��k�%fst�*8?26���'�Q��T���]*O0A�XC�����ctw&D�w~g���?�+nj% ���n Ж�f�G�m/�N"�������ŏ���V�(�T��g�t�)O�P�akK�[	Mt2���!U�0��|��jg�}�:KE��\=�{Q�tdRO�ؿ*tA��6�O�z�	�=��1j�%X�<7�v�D%������q�9������,�m�+�N�_�4���5-$���� ;�cv�i���'�c�ӕ�������J8�I����z�/)2��&{_w~:_k6������	0d�/�zO1�:�=z]��\Ye�'0X|����zߋp��|�H�Ll&<�2z������H�ګJ�x�u_\X���f�FД�b�Óg׫C�`����lV���|l�E�N2 !yp 7����c��&�����`!q�31�-X��s![��C�#�1<�M��Q���I��P���#�5��n���I�V�������(��nq_2�EP	�5,��C8,;q̳@�el����n�u& Ǌ�;H�B�K\a	�-�NUu��@�R���X�A����㫜�@�>�	6S`�	x�}~��̴�G{���»�6Nu��G�J@Ws15�1��;�2=�����E:��e�ب�� �,(��O�s쯗b�Y�qNٖ�ߣ����������g�>�WZ�����&w-3�Zr	I$�Oh�ͼ����$5�%F�ͅ�����cfi�Ry�U?^cE�����f1��O� 80��E��R[��VR���f?->�IZ�m�O�6\���ev	c�nIB���7ʀ��wU������O-��A�Y�iI�w��5U���s������9/����xci�����A���m���A[���ߟ�y���ZOč�Bߊ�u��מ���%8����[ݷ&�s�"��[,E ysD�%��c�sZ��*�@�/	��|�SU�@s!��T���_�X�Щ��5% �
�жQΤ���x�0&���Mo� r�����0�s��WN�G���x�)T�r�5, 1l�K��7o��
I����:�b����[�Su+��Q���`�ɠ�-\0�5��p1��-
�o����hB��\�Sb_E��LO�Gsw�=�	��⽿.�p0�3'�s�����ēn�m}UG��>0���ى�K���y�C	̢R�nD��D
������|�ˠ7[�4�$�D��3��}����������T�-��M�y$��=w� ���ԙ�M�i����7�}߽��V+�O��`,Kƞj%�G�j���*���)_��l�6��;���VL@�ǛK�V�M1Ncyۜk*��{cvc��.<: DX�#��^P�׼z2>Z��}�A�<�eK����Ik�-����45���K��C+8X��������?�8��_@�Zd\����<,x��_�a�zDx{�A=U7?:aB@��%N�"yM���U�~�M2+���L1{�W\��_gj�����A���$���W����ݎ�QT��f���9��ǌ�l0�� #}��L��r	�D� �Q����(o�%�Ρ
O��0��45�fT�c~�X\���Dd����1�G�T��S�haT[~��A�I�B�'����
����=LӕHВY�e��֔9"_�0��� H�yj�<���xi��_��ǌ�:�A�vo��o�;��]�x B���fq����bG��4�����7���wI�'�b�ф�J�#J𣼈y�E��h�&��6A�E�ru�0;�oc�$���?{����Ms��Ġ7v�� �(�:\��,�,c��7/L���c�G i�𜮸�4�C����]ھ��x��k�� �khM8Ģ\Q�i��|���J̱`n�>������rQ� ^�7w�J ~f/,>����+�i�t��,@�y�3� 9b�EbNn���Z-*�@6�!��,�j������{Sc��l�i��%=��ޟIP�.�ƀ�g�l-�c�s�"�N��;�#G:t��Uޙ"1f��n~���"�{4ģ���>C���y2k5��(�4�������c�Dn�u�`"�b��:��t���9��nf�W��
�LD��z�т̱��q��<�,�8�)¥{7�#;Yd����ËoO|�m�ڔ��x4AQ�!�����cHEg~�b1�s�T�\���-�W�f��l5]��h���vgf����to�N��J��1�l�c-��+	��W�;�q0�h�vľ9"V0#j�'�C��`p^�$6�pz%����G�؁��
���X"�z�iY~�Zn���y���)��oB�<��=ѻ�283������o�� Kc�l:[ �U2�ݻ?H�/�bj�x���ݬV����r1z+�mp$u3���N~� ���ỊE{�n^nF�\��:�R�;t����)HW �J���֬�l�J]ߴ���D[�ͬ�?k����p<�=6Xڱ���Y�����Se���@�T�\���a���l�&k��&��QG�)��w�z�7�G�'�_V�>yσ⩏J�աf�YO*	�Te�V��i��6���[?CKSy7Td�j|{�m�}�E|w�@ޘ��G��ZS����5?Zso��o�4�O��ia��ߘ�TF#���	�b��)aג��uF�q|�f��'��u����E2��%/�A���	�5,��3�@�)D�z&��z��2c�R݁} ��V������,� V@Q���K.|.�7=��$�W�4��Ԙ9��Ԟĥ����E����%����jJ�χy�"�gx� �]�[��T��#b�9�d��4^j�l��.\�c�)��#ÿ���IpW�����v�����~�j�Q[�'��ȧ��ma�z��Q�N�E�/�p˨4�7�x�8<촑O1}N�8�����,�=\�i��R�$h���~�4U�_]�/�7R�T���򷞭/�3f�e�Ʀ�S��14�x3�����7�cz�#T��R�p��4�ڑQ�v��Sh��1ؤ�ɉ����C��<~��~7]"�@�S\�_��zjg|*̭�kY|������HQ��SB��=��vn�0�̗66����I�/^�T�E���8�z��U�zy�cTj�gM�?��Jඳ��?:�t>P_t�o������t�iЭ]`����g���bH?#�Tp�0x=e��Kp���J�c����zJ]=F��x=�#�˺��ӏ�0�B�ʞJF_Q�~Wh7�N{��j�'��i�]M���u�=���'Y B%�;z�� p�6*P4���%`i8�[��A����b}/������-�ᘽ�5#R�Z�	#�sL��M?�U#�wӔ91�]�,�ƄtN�_�Q``yި�����5�6��J�_�F��.4�;�Њۥ�����0��r�z�+����{	}��m�vu	&?K�k�����W�׊��W��>j	D�gM%�WVU�r�������H���Q|�Ί�T�*�\��N\c|=���a�*�g���v�8�F�����BF#0�$�d�L�c��H:�/�@��a�neU��d���NTi�D�$��gd�˙��򆷴P�� n�Lܣ�O���=&!��)F]A�|D�!g��1�k��5���Y�B��hϴHU��Q��֯��������nQ�̋R7��n�(r�e��f�QC��YQ3GSj���W�7�~A2��l0QK����ĸ$�'��ge�R�s��7����&��T��مHF��	׭�9Ң���)|�*h�?��u��"�Kpț��m��B�k/��p��ѐW�EY�&w����j!Q��A����ۜ�K�bt�~�s��ڌ8�����	! Op���0F�T���WGg��/Q�Ү�s��ѰRb���s�RP�����M7I-&��x!7g��IwS��D��h[:�E}���]�{DO�"�wf:e�1���d����1Y��n��+����*�� CтG�����*�Y�Xdz�f��V��y�� �<W����YX#*(�:+$����͇�>�Ե�.����]tWh��([3�Q6�ybF�u�{����h{)�����r�'�����T;�������L.i��t�93����k7�ԡ�_	�gMw�>��41$��؄���0�������fp5���1�Ѻ;���`N}��Tw��E�r�޿^RI�/u���[�ih~��QUF�*E%:���ߍ����M���3򹭣�"���9��&��)�홂�ɓ�P��T�.���e+�za$1j6���
%��菾�U��Aؕ3�D���]��/�|6ܣ�#�I��\6k��1��R�T�םe��s/�ct��F�[��;k��✸�d��2��ݩ�����B%�5m�@��ɮbm�J���qVS�lb�G��Ͷ-#
t�0����&��x���t���F϶�����d`�A����p�1 �ܤ稧�����.jE��s����+�T��.C,
a� ���E�@���I�Z(F�H�0�,�Ҹ�����/�3�P&�L�rO_Oc��M�a����Ur�M��L�t�٭���`���������I�f��
�� �KIV�t�d��Ł��A61C[�1n���=�H��W�FZ�C�槆�w�z�^�@]Q5_�MU�w_;&�0GJhZ�<�{�h�0�'�tR�N-rkT5��A�p���#ּ��c���rp��g��w��#�V�/��IF:�ת��9&_��Ct$��]�8���7�aY�?��������#}B!��伆���ӕ߸K4�����U�#���8����_�yo�oA� �ځ2�~���B�-���1��6D�&�Ԯ|'��wr\���|�� QɁ:e�N�ܨ�@ư�� @@ݖ�g�-Ǘ���vԣ�xE�ydxI��!�G	�����۹�P��)���Ԩ-!�@�S�㉚�)s1���x�b�[�5����'8%4�zRb��, �F�N"`P�Q�Z����
������K�|���F����PfkP�g����t&S}ࠗ኏���O�97��!k��kځH��űD���1°@;���q\�|��Ó޾��\�M�S�0	U����U�M�c^���
t/�(@�/F�4]��s�A�j���7�I�6>3�s�O0*wDDЃn�������a
��7�!��i�Tƭ���&�\O�x6�,��I�\T�����?-8cd.a$�|w��n<�:F�޼�
Vͯ �Np��A���b�S�c�b{��L�PD1b�dU��D3�}W���j�9Q��s-?��16 �oq�a�Ό��,�N�X�S�_o����rص���*�W�}o<�/��u��I���j��c%N�`�>^�@��izG{`WG�mT�$�a$[QҜ=k�>�n&N�����dc���L��=�gg����aWA�?z��U��C�dx�e�NB�`|qz�g����@G�1n(u��������^4��>�t�^އ�_ 3�4�HB�{��F�«W�e$W���~ګ�ɣu,P�Q��8��.����]�"����,�;� ˮ��cv1Ĕ+z�P�:��5�AD���N��0@m�0��"֫>O������A/�z�������~��Uw�m_����9q����� h[N���3Y�nA��"�|������Y�?', ����3�����L�ףٗo� �7���+-o��*W��;�\��+v���|��K[�\�T�ݺ����]�6i;�X秕���/��y`fAF���!�͍�KEʜdV�T[mP�/��l/�������U���(*I�����j>� ��f�!v7(��̰���_����Iޛw���u��T����iu
vG�������n�1/�D��䁚2���r�Eh"�ˉ�Ӱ}����
	����k���pgL�7A��K�q�	��F�U���$����!�������wp}+G�Vj��2 RԀ���5����pI��J�:V�t��0��} ��\�r#��(r�����h�]��/m�J�N����F����WM��S�5��1�_��2z+N����k��;|Vc����*lp��֊�U@x���9tD�OS�5y��IgO��6�������f�т����	�� 5���7;��&���^�����7k����)�p{�$K��ʋ[��g�+�.����H2�I�{0fv�M�� Ub�t�~_�&��T��w늇���b.�(9��2" 6	`��W�o+��Dz6�����TӠm��ʌ ���o����v�c_�s�"�%�?�D�OdOV��f'W˧z<�D��O6�Q�M	�YE	Ὀs���G�qs#ُ�bq������);���4�M�%}SG�cٮ"��nb-6e��G��/�j��nm[���i�<\�?�����T@�#��|)���)@�E�%�x�ղdw��-�g��8�9bQ=�05�l~�a*�0
�=�E����1e_�R�.H>�IWZ`o!٥Y#�����&]�kl1�q��cc�Y�WT���}pS���k�k��}�2E���EtLg��2Crk�F��85JN���a:y�CKɰ�zm
=M���
D��o�X���N����~n��hhO1��DN��S��Ex9
�&o�b��sK��j��d��(���mxE-�NLX�'�M�z���;�����Ti�E��
��=�B! Q���<���|���<������n(��Xe�ǌe��2�
_w���H�$F#�)z,�T��*sӫE��y��Cs���r����h����ե3fq��Y4�# ��01]���^�5��]�+�[b�̋﫰} Σ�o�,��z��2�[)�Ћ�}�9$W��������;g�HK�*�GM�:.~�?D���Ek��#�e��e�Ї�ǁ,y�#�q΅��������_��.W��!;&w���3�yo���<k����z@P���r�レ4���T�8�5Y7�1ǜ{��CL���^�j� )V�#��J�h���e:�\�q�<L�u!�e�;k
0��߷���h�P(�=[eS��-4J�*B=�����06������}�xŜ�U�6�"� ��6l���(��Q�m����pz����%:�d�ώvh8�6�d�:�z�Šcx��kL$��]z�~����V�)n�M��<x�� �YA�Xd��Vw�Κ��p��89%�a�l�l����`�3O���;���k3�'�m���a^Z8f[�
��X�q�]��+@G��C�
	���/����k���@!w�IF�� ��uƎ�a�^k��-�fԝ���zR˙����U{{��?ȿG�!RN�TD���0��Ū� ���ksW�(1s��0��S�3]w
�6���)�ЍR�</" �!� ��!��O>z� �qip���� ��/kcFK�J���#;ƇE�N&қɠO	:^*���j9����U�1�vg���oCZ�a���􋻊��}�
�	S$q�j{�0��۶�9�����;�j�IT�K�z�s&�L���x��U�`Bꂹ����k=#[�ɵ�� �s�#����8���AT���r-�#n>���܄m����E�K�H���S�ɠ�ʎ���wo��ψ�3�ġ1¼h�e�O����`�H��\�b�7� s� �}PfUut�XG4�M�U|�9���Û髁ނ��S�~pJ�1meK����Ҧ0�Z���=�-Δ*Y�[��aw����