��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C��(b�g L�N�W/u�b|���@Aw�_��5����w��&�T�`x��i�>+�_^�u����V��0�d]����w�������x5?�\.�r�A�O�R�s��H�2�z/�W}��\]�����8PZ���L=����".A)	H���/���g���GN�����G	BX	�f����Je�|��t�!���s?.Fݮ�Z�_�6��hx�w��[?�z�(�7E��n�7������8��M�g��< �HI��oߐ�9Y!��!;��@�sy7�g�}�o����'V�C'� i�,�����M�8�͟Eo��_Lr��s8|%���w����w�������P�̸�	Ȓ@�E�B���a��Q�qwJ��k�ҍEүb��u��	Q2�t¥`i^%/��2|�)'$��_�E��AQ�/�*��^��E��#D��e�v����Q��3�u8S�.g��u�\����#� �@���}/��xW%�ᅩ�f���d���W��W�L���'�#�O�9!�f���Xm/N���O�]��ZMD�r�y�i��>��B�^�F��}��7%t;uJ��_!ap���J9X��tX�4a""��g[!  ����C���U�J"H�Gn�s��OO&�(��,���'}u2�<�2��؁@D�� /���|ꦆT�,G�9�xrKPQ��^�*~GʮoF��,���]�i.�������wDK�$�ReOؘ>E�$~���V"-����q��������qzS�¤�f�hTX���u]K��C��-?��Kj@���� �{g0����lN;��,~�<8^�5�P�҄3���2�(��7��^������`0~s� �%sn�M$�[�R0-��Ừ�D"MF$��V��((�d�d��^��sԕ��˓Qw���	��� (��oы�E�b�;�
�Cgv�Tv��V!�\�O�K�̮]�����Z�ڸ��hdoɵ�QkE�2^�����4vD�p��3�'�zm��VB`��5(ʍJ�ɣ*�V	�W�����̆f���ڪ%Pzg��`l!�c�����Ky��?��G�c	dg���%�>���|p~tT �\��iz�?�k�__u��jh7Ԅ(����h��);��|��SS��S��br���P�J@��.f]�ߝO�%�	
ۜY@�,��U�Q��<����Q�Z������]�Ū�;�o��V{\�o9+�VB�W/����%�$Y���@\
{NʒL�Pp���������,�0�.��).��B��ɕ1F��h��lC��bn~�Ѿ!}�mC}>2�@�^+݃}��3�1��V��3a��y"�D��->Ŝy+��c\�ǋ�[��x<�M���c�����ߙ�M���9�w��n�˝u�=r�f1���'��V�$M5Z�kGN���Ϛ���I!8<��Ϣ��	ҷ=��IH�$=���)��@z_"����dm� �*��\F�5��,B�[�`)d��A�C⢊�ɍ�}�e�y*d���+Q�8iWN�Ǩ�U6�"�2N�+��+WU��[��5a��H掋��S�"Ņ��t�&v8�rBM��wr�Gq�����H�-5�A�6�z�&���'������g�Ξ��?����4s]
jf�^��>&r���K�����z��oҒ�Yb���Μ`�E���KCq,��l�BK��~DG?��"D�#�!�$"�� � ��2��O.)��=��6a�U:�F>��N䮂�s����6��<�'�w��y=�g��.#��Ytv� u���53�B8ǖFAj�7����F<6Y��/�tCĨ�3�v�_3��Y��Sτ.WBb�S�CYR�|fZ,-]4-Y�|owC���m���A֌6,Y���� ��G�jH�JS��\(wݝ,�@~�����pmS�b�3��Eq*9	zO���Q_�X�;�
1g6�@�8a �//G�A8��9.�Ჵ$��@M�O8R\�3ŐfMA���Db}��4� ��ir	\޴�ӵ�)~� t�����!�崵��h��P�V�z�kL
����釺P{�7٭�.�D���`�Wc8�F��O�λ��n�����'j�2Y��5<�5M&`vZ��_:�7
�(�)ڀ!�#r���4�y�}�/��7n�5�M5j2!-�sr��O��>����ri�E��7�����@Rr�!�)*�g�&��d�}K��bǝ1�5�}dc���f���@�R/�|O~U����R-�h�_�}��mK�h��>vZ���¼Z�8g 5��E(z#�Q�7o�'H��8��Er��!-[9 �=����pS־���[��Z�e��u�����ó������p�%9%���dB��%i���X���*�Fo�����\,�~�Ai57b���6#��a����~�&�K�%!��\E�j'���ٞ��kf��������a/bL7�BU@�;l�4��{���.�&w�+�h�j��Υ�c�PV�QN%F��d�nu-~i�mX�F����0�`$��׉�32�u�pO^)������ +��Uc҃�*�a�bZ��������0uq)�Ob$�w�Hb�dn
�3��E\�rV&o9�m�U��v�}/���"!�����?�f��=.-��rG4�m	�MZw��+��fZh�S�/�ԓ�ܽ�l�M�$�@�q5y�;�S�x��z�=��΅�5�Y9���`�=W���K� ,״��}����mU-Kn�����#{�+f���U{���IeE�~l�Yݬ���m�x�gb@���°��%Cu7W�iat����p��'s�.,_^�X��J�����T�X�G$���.
\��톎5��!m��ˏ<��q�Hچa|� �K�<{�°v�T�C!��M�>������_:�鿲pS%e1]�&~+��H����iJ�Cr��*�۾���
(��[r_�=y���(r��.\����4UIRr����C"}c�����3%��ED���G��n~H9��?�G��zC}�#�<	��*?��]�?�r�8�L��\�_+A���9�טs�s�Xkh�����g3�I�V	5,Y���s��J-���z�UC΄�4��ȁ�jaS�����{[Z޲��!N�\��Ũ����u*;����$h�%�W�steas5���~Od%�&�u�e��?�Mac<��j܏Qo\���/�]\o����`X�s���sY0\�ZT��\�:Tt��{i\�ϔN���⢆5|.��Q[#<8��X��)�	=D��d��(�)�k���ُ����/;p����e�PY�F�3�Y��̸�c�`;C�ұ�zT�@Y�W���W��"�f��l�H|�aA��K'�O���$FVr�}j�7z|Y8wr�E*��+8z�kf�֫��O�(�o�ΰ��^AE%�V�w�~>3�Q���i�+}$��I�.L��tq�/1)��e1Л���6*��j�G����f�`3���!K��x/��ޗ�N@�+].~�e��X{�-^R��J'�~ߣ���ݗ�#��3�h��t����3(��}��0e$-���S���?�+�Qط�b��|�ՒP<�n�k}
Z������ʳ���-@�q�[��Ҿ}��Y�7nab�!}�B�_yA��x��e�1 $��i����/��~y� ��QhUjGx!N�c��J��%�Y�%��*|4&"{h7�ۊ�~�;>�-����Ţ B�=���r�I|sK.f��0g��k����4�/��N����A�����*�hGW��v�w���<-b�ٗx1�7O/n������ tC���m��cu��|�����k�Wᠢ��b�t�>z�Q��u�$9d���L2�d�����w�܅�c=��BR�1�Jv\$�+7���]s�꓎���"��ϦeL������'y���f_��jd�!z~͓#������ZK���+=<9P��(��@��[e8��;����i���F@$��^"!>b�dB���s��D�.^K"�L�@���!�z���/�q�j��n��v7K�2�g�5J�
�V*���'�s��)�P�.�;e1˩��D>�ڀu)��3��Ih�<�@~+�� ��1|�$\I�i����y#��e>y{6�Hu�����49���MJ#�kg�s`fJV����5`�SؐC'*3`so�Q�\JC�['�y�a������ү���,���	�G�!@*���!m�^b�e3�a�_�:%x\g(ݟֈV�`Q/C��Ze�U�><� ���b`+�6��f\���%�\��_�
�y/N4�N��xL$*
C��{g�-��)��_m�
����)uKS�F#��_o�����Ja����G ����������<0U�J�fMx�~0�ނ�����n���#�gq�ݜ/�����1T����n��4�;�#"�SU��K�mM�"�4���ǈ9�C�t���}{�� D�k� ����bj�sN5S�]���{���`r?d�L���us������&\`֩BW��uE���d�e��|�/ު���{\(���zP�3UQ�r�|�h�x+%��4��|��p*��[]gR�����$��Z)��!���)��Χ_�a-Xd]5��S��Vq�l�M	�9�HHأVmS�(�{v3^�h� �;i����-؈�/�;���=4`g$C�Fi�̷�w
���8~sc�A���K��]�0��8g$�����>F��و��y�,��mA��SZ�=t�҈���Jl7�±���ù{-��հg����T-m����qk�2T������Hy�	$��c��K����0��~}Y	�������vB���]�^xŰ�BG�����5|����>vB)��R�Vby���|�[����� m��<�9_|���0���B����Φ}ۛ|�ʴ̈�rp�1�w�����F�e�Bi �,�.*p�]�z��F��3hz݈C���[�_��}�� /P�Р�bϯ�]�Zȩe6�H'��n ���T�`dCG���s
�˸�=�/�� 	)��><�1�ȴ����Ȥ�n�U}ńS\P�X�Y�ڧ��M�	+zN�&}=�c�/ݴ���3�0��v�&-M�@{t/�J֋� ��RA�F&���]�P��D�D��tyX�>��O�n�+��R�}��m���hd٪�Y-�P��|�P
�C7����#���g�Ja�M��"�\Ϭ�L�U D����t����ZlJ*�A����=q����� n�H�V7�	�.
��m�@U���b��ɤ��x��7B7�΀���,���A>�s�:5��-����y��4�7Zh�
8O��xg/Ù���W�#�R�~��]wIיu7H�V%�1����B�!&���A޾x�M �6��~��<�M��8�d�ܿ�ξ��K]����|'��uŽ��xV@�Z������dJ�����B6w�<6Z �iDV�\V����X!�R����#�J�Aj�Z"��	� G���PǗ�mk� ]�_i��`�L��
�l�P�Ja{�wt�qg�3�P�:$g<G$���#�Wiy��F�\!���2����$�h��{���~s�;r�4�:���P�Z�3���\G$pd�,�����<��'~B,��jp/��qf�0���6�3����u	#�3�x�Xs>�l��sm���g���~��j����U��0b
�wY}�s=�o�C �W���oνG.G�hJE��<Yq��޲��x[�G�-�&T�x��\�Ql�\��i�����/�^�*n,w�Iu|�]�ς�/�������N�n���Ҩ"�	��b�Ek�'v��T]��g�Dr��ml�co��/��Hs�F�O�D6��TcHy��_�{ޭ� ֐�>y:�lW��;�|9���:���&����u��M��paޏ/��3̴WH9<�C�L�]J���6/�=y�a؃{�K���F#�vZrq��@ҏ8o{�2��ci�BC�E8�����($��
 �n��r�
6���9��	�;~GG6�+��-�	c�G��F��[w��@sd�b'�w^&z���ҿIympīB��6��_�����!@�3W�3<Yː=O�XY�Ɠ�������k�A��CX�ʍ�z�[!bRO:��t9J�/m�ɑ�ώT+Z�&8����F&(��DMx�e��[�3�%f-��Bl)T����u�4q譅!�\R%���TS���N�&�D#Fe��" ��$a�N��XGϱz���F��/�y�!3�[��1y�� �E������2��x�U��31�1>e�A|�\���E�i�HnGCB7�C��9\bKʖ�k�����E��<4�h_����kH\�sk��q�O�� X�J����FJ��z�.����KN�>,Z5��m��c�޽�Ժ$\CIh� �y5L��զ��a����(����Վ��M'�5v�7��:Y���5�~�p���:P��B
fT�cOa�X �m���j����&E���L��i�\x�<���[�rY��8�8+�si0�A�N$M=�"p�y��{��Y=�P�$�܈��)��{��}`�@�	�D��o<�{hA��BD&�yCe�-�0󃙣�Ro�n����hA?~D�BS ���Fb�5i��xH�t6��C��2��O��+�sFp�X�ȉƀ��-׃
�ofp�37%v��*	�N�n(���DuBf-^��Ĭ�K?A�����P�Vy�`�S� ��]�_x���B��6���t��22����\0�+8)ݯy�<��qD+�����^�7acH$΍#I��c�
<���S>̪��2�f<�H�d��4#)�
k�v�/��K<����U:�`�k��?�ō�V����x�=MS��ͩ�z��'�G75�EO�.�DkY�;u��s�RO�C5�n�vKA��^w�wiM�� ޥ� ��-/��W��~�;O�z?No�����d�=�ֹz��2ړ�7wAA��72��*��Zy�H���k��a?����hiJ��pZk��ޤ�-��y(���r#�d���P4D:����S���u�a��Pحqeb;Fn>F����@	�Jy�M�����4��u���qk
�Y�Ѳ\DŐ!�ƥ�c'Ϧ��[v�ʂ!i�
����Sp�i��ʖ_��o�����a�h�`{��N���ON���Y�i?-h�.7�u�t�����AyR/�	R�UN�t�z��8+�D��{�s>����B��ż������D���Eҽ+&s�swQd�e�z�o
�.�"�^�߽$Aݫ� H��mSgs��`_U�,x�T\�s�SVhLM�E������|x]dZ�5%-��uGO���_qb}��1ؼ��%�>���#��zA�vD,�oq�QB�^��De�F�QM�&�HE���4�#Lp/.ir��!�ۛK'���to��K���h�t[�OV���Iߖh0|>QH/���ǟ9ZoS
r}�����[��C����^(|89���k��F>=���� ,9�VC s��7΄L�/���Z$O�\��kWU��֯%@����*��z{_���Õj�D]�zJ�R�쥆�V�D�<�G���^�v.珁R�$�RQ�+�?
b�o�����;Sr��ыA�D�SEV�ǜ���Ҩ��9J�'�h.3;}Q3�B{&�5�%�
bI��
g�o��Wo)ʇ=�F)��3x�����T��oJ�`�?�yL�o���=@&�|/�5a< ن��B�,e܀꯽��4�pԂ�H�/�mw�dʒ�58Ց��Jv����x������B{�(˨�)y�t���nD��m�8A ����}޹���V�-���N�c���1t$\�����KՇ�6��/k���1l�O䀸߷�J#�;-2s��*���8�t�gE󌵴�-W���ñx�G�^o ���6q*{��1%L�E��������K�Q������]�3H���y� *���d���gA�F�5�c�oz��Xb1���KG�_B����D�=Q�R�4�;�giCX��6{]��鹏�|�#�(j�%rYsr�Ѽ���h�]��4m��,���?��U!@�W��ʦj�#�1ڋ�C .�\�%p��~�T����b `�p^��Ph�F�y��+A�ۀ_��O}TC�	D�5�:� b��;s�[`q�tjo7�x��څ2s��>Ki��1��D�Ʃ��@~��9�_�����x�(�c�vtU�m�ח5%U�.��V���>pR�=�W���s�Z��[ �-�.���]�±E6\�x�9�#�dT����H�e �<d�['3��7or��_{/A&�kp�L��%�+���ߴ˗E%��.ɭ�g��IY�S��Q-,�~��pu,b�3ŀrc�e�Mw�R&kƜw0��w�T��`J����۴��2�4m@:�2��x��T�ij�GH�(j�\��Q��GO|�"�/[l>+m��J�An�	3��|�z����ڴ?m����f�Y�q��]�2��VtJtsQ~�2O^�ĖHa
�BIX��⺩��7K��4_�l����N vQ[f���H�r��|l?;����=i�G��5QQ$-�Ű_��1Q��&��uT�^!~+�%=�rN���`|�P���� ���}8�e�D�󵫜�]��T��nm������N�v��Osfo��S� yO�J� �)9x%M�m�5{�DD)N�$������wo�wDɌ�,@N�w�ݩG/	�� o��\��ZЀ�+?Ot�8ާ�Ax�^�ck@���m'��)��Ia��=,%ܗ��K(��橧��7���x�P^��a2�畻񬴁F�@)>�JG���ɔ$1@�����٭f�n �� ����@O�cЙld��OՎl���)� �� _>mh�wa������O�o��5�Ҿ Y-�?P�9������,�}P,�x��8WXl�`�섛�g����J�E���t�g�JS� њ�0�}B�]�"/g�?�UW���ַ�U�(���G��|�����Qn��;4����p�{f'��,�w'�A1�Q������
 
i!���8� ���8�no)��m���J�>�=�G�S�ʴ�ؠץ�a�u4h.OZ Dȏ:�Kjk�1S[�-#[�N�;/���[n�a����0�ҧ�,q{����NM�ʮG���$�V��Z�`���x4=��<,���7��M�	�A�_�'=I�!��2lZ�m.[-����n	�3�1�eO=9ah��1�^�!�SJ�n��*�)=��'b����3����s��ff�G+�����q��ۘ�n���Z�Tx%|xT!�Z��<YwBO�ƚ��h{����q�>�P�l%�cP����#ٰ��Y�� ��\�I�Q�ኜ�,���-�T!s�����Ӻw}��4��A��M|�Q�n9vLڿ�ax�uƪ�tR��<{��*��ǿ���/��ު}���[N�lE���(��r�����ίQ6�H����q��aE�a��9 ���(s�Q%O�@F���l�m���pݒ�]�1�roK��{Ǡ?��z�P^�YF�'^���� X�� M�{<I���!&2�����Y�J_��-��L]'��ý� ��%�!��!=���v�W�%k9��V�������f��GK����fֿ�&��9$�����2^�'�U=S~!�	r.��ͦˢj�NWTPa]d��m��UP=�9��җ�TT�%�}k#� y�/�����v!�u�Ӆ<*왲�&x��R������=����:��0Gu؛��L�����zƼ/*7�~��+�̭����b!H"@�X�۩y��.���������%�w������lP�g�7sh�����O�J�s��+rF��x���N��\zD|d�2|���7��������#y��7�����Ed���c;.C�"�l��T*��[3ˉ��Z1l@���	+��hW��~��
�:����u���W;D �;�,o���w2��q�������?�񇺋r-��Z�_m�~���W/�%���$�7����|�E*@�A��y���Ғ�I]ky0W���񏞃3�]�+�6�I3��0���V2<�Be"-�c�/>���'lI���?�+vYl�و��4���R����q��:��`'0�!�Z�v�YK�r��ӽ��T}����vXbdMM����3��*����_��Ň��R��j��>���@&�O�yf a`[~-�CLE�U��~z4J���J��k���S��V�5�1|? m���つ���hǿ�{�Ep�U�Ƞv�Pay/�q(��~R.������>�\�W�{�|�(
s�NB�܇`�Y
KS^�|�q��K#*�����H�����~����o4lV�.���ԃ2H��SE�.o1��C1��ѵDHA��85�1�߾4KE��!�(^�^�	��]Ϩ9��H���2j:xp�^�d|��8s���j3���@���!&��O�o0T��f����K$�VM˶�2���\ԃ�Q�w�RE"E&�a���Y҉	 *��6{�2�:��I��z��d�)��Du�=��5��0#+�5	5�s�1Q�q�_���(�"�Iӊ�|�C6����?3sE���PX�XRo�����-ɶ�)m�@$��1�">�/ȁ�Rֵ����CS��ݏ���J���f::ehDBP�r.����޶Q��<��C���M�����!�A�������hs��&���b�
��c�\�ղ+Mא��(�gd�Z?׼����I�rM(�@Hdp�\�U��[!�1�)�e��n���u��&#�bt�C�Iz�@���m>�	�~����^�˷!f��&<�,�H%̒U�wp�
˖�O�գ����
�<��7�Z7$ο!j�tжO#�f���������(J�����ʫ�,���w��,�Z�(���Ě�y��R��ǋ�O�:q�|8/T��G{+�9�����й���;��|�9$<�)��#&�6�^)@hs�\�߉�YhgǍ���{��B��W>X����.	S���h��-���FR;�w^���+����
[S�e�	du��A�d�?!��mbб�$�}��wy�TA�&��Uj�=��۶�X�x�B�Y/L���"��xplU�/=�E,%^ԁ"�f�[��V�&S�q��*�&���fJ/%0L��w�w�����.��(�G�L��M:yo���ؠS9k�D���9��|f8Ѵu?p�Ӱ��.h�PB��Qc�l�����[�ʧ]�!�i�@��	ؤU�Q�=����I;���#������ط���(� �����AO�}��K�^����:���D��x��Iݝ?zĞ��<�߆5��Fo�xc#�O��kT�0��#��pmx�k�.�;S	����'�V/;�c��հz�2a�s�IcѪ�g,gz��K���!�,@�������� u{��h���%麐B�z}\*
f�k�w��Rϡ��+�64��-5`���|Y�10��j����x(e���'�����I�j��J���7�R�!z�-���U� R��X�d��ʪ��J.�v�L�g4�v�{��Ve�
��� 2m4����CK�{�*�׼���<2?��s����7��^7�QY��o��J=�n�k�K��ɴ�&i�1P~_�'d,�Iy�Vj\S������X	��Oj��;cᖔ6���5�������1�@����VG��d=��H�$2���|o�#�?�=f�#�31�a��#5�sL+�������?A�N,�
H����h���v�~�}��#�G)�E�4vC�v� 5or�rC&a�7�y&�����0jy4�kN}ԏ�F`��	��jǛF�Q�$p}�*T������(-��l�K[U��Q	�)+�P���j%`q#8}�qp}\f���[����n2�kՎ\A!�xE>Q�K�z<]&���!�W����gI�;8�7��ЕKɘAx��h�0O<
K^��Ռ禠���BJ�3���"*Y��:����q݃jN�_IfN�$�"��(��S?��2F�Or�@`�Bx�EASFA�������ʓ���h�R��H��}=�wA�ҭ�/����