��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V��wg��+��1�0��"װ��_�����/$j\�4�eWL}�:�Ԕ��P���	Ȉ�P.#�/;�b����j;li��(�(�^n� ��q&�w����+�a���\��J ?#�r�xtܩ��3�}F(P��G�2�H�r5�$�2FQK��@���I\�������ސ͇�,�-�'"U��b�'�(	�s����C-dO#[H��.�N��|�9�>���sĐn��K�A��?N�������Y�j��3�0�!��߽�p�a�7��D�a��Q*c�B�(Ӣ�K҈�7��wB[�U������Gz���\\I�Fܩl�0R�T��-c�
�A+�K��j��FD�E�82ǣ��}�a��IM����lZH�am���׹�D룺�Q�9�6�g�(�p/}J���y�eV�u���\1<˛ʤB�+[v\a��t�_�Wե��g^cu�����R0D�R۽���6�D0R#4`�����_���8�٤(ߟe@�b��K��o~�t*�0H���7�ġ��9-D�e����3#�'��?�����'9a�'<����R8t6�U�}�:{�s�� ��p�[�n@�(^���s��|hr�&�kv�Jv�h#
+u� �d�>\�
U#�H�c�3c/�����^c��kO���􋁹�O=��6fw9���X�ˀ���3F����尗Ư�]\�$7�K��$WR����'�8D`t-�C�*)C� <��x̫,��_�
�9��Шq��qA�
R�eOB#�U�e?�Oҹ)�U�i)��#�Ʊ���K�6�Mr�4�>����5�#D��?��Z	P5�W�8��u��L��#��.&�u�(L@K�L����zο>f8�cq���W������n�{�X��;�Kv=�"��di;�n+�Ѕ�5d�F�I���,�iB-�|��[�\��C��1�R�ܴ�Y1%��RNdN�`�4`}^X1G��}�X�8�U�Ή؉wj��!� �kU�&׋�W�I�/���9*�� ���(���1z/q�<�--P�~��Y�r�?Q_���k�����r�X<���ϧi��L�5�Ư�8%�v#yG�9� �O�	��㟾��G'
�d�����e1�od�F�&�ϗ�eqI��S pa�uU#tO�~3���T���>�b�%Y�&]�Ց�G��5hf.�]:T�]��iQ�*!�o�x�c��6�Ԙ�aXL{�-���V������r�bhD����7�������q|�vl
r[Q|ƒ��`�*�S+�*��8aT��G ��K!z���BU&�"�tWB�a9�h�fT7BZ�����0�E6��t��`���*��YV�w�̫]U�'��!�6�;(�G����?:S��P��φq��[Ȳ1�tV2KI{��Mylo�:��U"�RѼm�qBWH�B.��,d&Ⱥ��A,"���X�"IcXiPn*���T��aZ��{eM���"��I�_S�-KX��!�,٠qE��b�XK��W��c�C�L�Pzx&�(�-�������(��Ki�p�������d,��4RC������?R���|?���	�`�~�8�7�	��[%�Ћgm�b<�oP*<�xwm��f��->�|���L�2���0n��	Ea��?ٟ�.�%H�#m§��@A��\�Geo�jؔc�
:��O}��)��p�I&���y��/�k޶Ǆ*��v�KK�ZAW7o��N�������<|���1e�d	��N�!O,��9�R�؟v�������ئE��ND �W%��� ��c�1�2"�2�}I�1֬�
Z�Rx0�{��]aIsZ4%�4�ңO��@Hc)D�t+-<,���k�
A
����Y���U��ٮmR��vL�Oy��/��a�q���K��y������ K%�#�2���57󤛥���p|�6R�f��������v�a@�?_f}1���/�ӌ��]�h/�7|�	۹ X7<PJ�v1���ޭ1Wxoˤ'pݹ&�i�=���wΟA�]�{�Kr�!;�cr|0^B��]զ,k'5}&w%�j�e�?ׯ����s�tS�v�1��o30G����҂�,2���<��*
�&Q��f���6U�]r0�����SE0�y�.9]ph[�"V���,j�"eh[��,յo��m
��iգ���B8��s��zn|��P^y����f��̱&����[�7��
M&��)#�b�������KF%PP�G�v�����X����O�������60�M��-h�Ẍ���I�0ւpB�MHv���������������z�D!Ъav�+^����J# ������ށ�W@=��k�%�GA�#ɖ�ӖM�ٖo�5�-�̴�@R������^5�yDi6��3��PɑN�����T���E�3�nnmo�o�O� ��щ���uy=�B��P1���m�����ʀR|W�&��Xھ!eŏ���:c-fg�q�G�<�XGetP�r���o�۷K}7��rK��i)�R^�(�����§��m��B��>ݖ	ߦ��`ׯs��ڔ��>s�ߥ�-�(A:l.#���X��X�nS ��zH�������[�+�8әp:��IfI.��&�(Jݫ������ac��/H
�N~��R}d3���f�o2߶�Q��n>5@CHR�Z�v*0��s���sR�:�	.�n�)G2�?T3oBC��H�@�O�O�缃����=j�΢%u���h�+Ht
L,e=sQ��<d�
������u<u��vuo���ƕd�m:�1�8��9�ҜoMh�m/�o0�\A��s�3�&x���&M6&~<�9������u]:��Bt��4Q�#N\Q��Y��Ry�(��O2"���8����o<xnE]l$*y�������R�9�hFf��3��3�����GGMP���#�E�J��lA͟�[����� ����?��b��O���	�|��5C�W�8�wf���=�/6��r�;�D�1��݆p�Qѡ��x�4kI�Qش�P:C���BL�0v���u�(�Z\�d%�)ʻ�V-�gF��D"��:n5�!Y��n���}�9̅�R �@>^����w����M�5��}"�1=u�C�N+��V�q�v�\X���*i���G�8tKX����&B�m0N��s�ȳ�ߛ�,}?����:��)�&n��Ǜ��?4��.쮓���j�W�a$��(�$�w�����f��?�MpA� �����$�Ƞ�m��4������V� �n�U�#lL�8sE�;���Pi�d��%Vs����D����\j�f�ә ���L+�Ǭ�