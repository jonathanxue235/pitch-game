��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V����hN=��a���)�硹<H��׮��`̼��D�g�;�mR�#rj��S��k@'�q�/�ha��pc�R�(��g�F�ו�����`d%D��G�qK�DW�+X���iv�O�O����9�t�0���`�<�F�2MGJ�g_Ю3����Na/��4-^}��ru1������>�9��& c�dN���(�lE#�)�<�A[z�z���rpRر�ɏ���Qdɶn�Dx��jB�Z�}�0���=t�xx^�����O%��E�l�Y��X`�24GU����W�VOt\�5�O{����fw��+�+�� x��Gv���'�_��}n��]���g]���2�sJ9`&�� 4SǢ��6�S��~2��8����z:�Z�O�&W���G� 9��(t��$���z�hL��Cm-idϹ>�u�띇�;���JIE"�~fO�-��@|��.�c��͎�ґk��B�Y2�a� 5���jcA�3�pޏ凰�D��̄cdh����!��$ ��e�OF�q��T?\�M����08_5^p�o\iT�� ��{d?��F�pV)�C�^��,����SFJ2PDg��.�BT�5oWU��o�`@�N�SԷ$<�=��;0�"a5����_D/�jᚩ�}��dˆ)p�5*�L��`YF�T5���u�^v� ]XE3<�5V�6��%1#$���J��<מ��G��{7C�S���l`���-G�j�r.��t_��h���<r�̀�� ���ku�X��%�D��x�,&�o@��Mm�~���7�4���I�W�i��tN�0��U�W���(|Iyd�a,���D��7E�2A�U���� b)5����&�kY����U��<nv��O>p��<�lb?���#���lK&�o��W��j4�Xrޙ���Gz�O���]b�&B-1�_�7lW�U���u�Ǩ�2���}@�>��r�	qɪ�j��N}n}5����� x�<�\�^\�(bIt�ݻ�8ꡓiu�a*$J�v(���t�ל� C(&L��Y�7�lI��ɳ&a�"�/����m��OCqb����{����_��+}G��˸B����oA��3_�R3VxK%Y��-yc��)E�������z�RsqV3��.��&B���\�$�s�
��Z"�{��t�\����>E8i�l�;�����.������>�?�=��:4p��}�	�
#ES����u__�򫢾�kd��� �����2l	}'L~��X�ҏ�s��C/h� ]���a�(�ਯ��>[��~'���&M� :&���:u{����R?QprL���/�W5-1Z��>l�*�j���}(�{�_T���ɨң�*1o��H�L���d6�n�ʹ�_���6W܋��4�+i�P���[T0�g���)k�䱙S��0�¬Q��)S�ol��!�h8m�o�K��~��pӲ���(��c,#U �鈠b��f��j�j��x-ݼ����yU{���l�� ^�w(#QlR���T�?_�o�甀�)��|��v���I�D )'x��`�m�=t[Um����c�W��{��@��p�
�'/7�zkQaÁ��2%���(�.$�o�+2��E�V���#�� A���&��Z?�5�]��]�GJ>د��*�USp�9V���-H#�p/���6�:���f�bK�8b��ͩ���B�RKi
_���)����=# ��]�w���4�>�8�e˄��k��8V���A�t@Z�T��Ą�N9�U�K���I�� N�ۚ�d�� ��!�ɘ�'��ݦ��d_�}[�{�����	!�6kO����m���`��y��ZJ9�+���\-��VM��~� ��т�c�NԱ�S��J�"x�5?
���T�g�ar�Vx����[`G��� zV(����U1����CWs��@4�q��9�l4��<���w��~��((t�I�>p6���햯��3
$a�]c+#�J�>��58F���?qS�RFK<��9�Ѡ�6it��DS·�~*-
���L����u6����#���{�,'�J�w?vPǱ�ul���x�>z�nꃁi���ڭ㌌�(�e�6�MY����P�G�͌���DuRZ��݈�<���8U�^���W��}o��q��M�C|Dlpj鯾�>��^N[M��+�7ҧ�&�8Q�x�ZCGϼ��Z4u�t���ܤ�EBe�YKD���1�l�xaRnZӿ\,�*\Js�L�X)�1�N�=vތTb�Zem��Mk��\�&�7�b;13b&a����<tݜ��Ϲ��Տ�4���~e��:ͩz���gn9�n�j嗤I�o���]� d�<ZS�V�N�Qj��ͥ?	o�V[���G�pA������5MK���#�p)����*6���c�6 #Ŋ7o���O�`�@4�on���P4�{����~�ɡ��~���+"s����.�*���:8�6˘���sx�ɲ_\7�(5�k�YE%��ƉD��P�-$t�DR�i���[�4��sVi��V�ֻ��c�_�a��s8_8@�DU����>-�u~�o(ab߸�;��{��O��Z�o�� �a5w�&<���pWm>�HH �d���5��=���s�C�J������n��'�_���KV��Y���By�w��m����g���O�w���T��	���r�/� O���Cz0�H�<��@��$`\�to����4z�sʒl��{:�l�C���T�e�T��@��Dh<�M��L�ԖלZ��|�:��m7�����c �%��|�q;o&�w*`�2!��Vrr;�~��t��t�=nݽί�ŭl�&��^����p���l�����-�_+�*L��0�faM���C��W;j+95��O�bՅ�;�G�>篘f��+j�f�=�:�O]M���Ym:MEc�C�#�.؟(��2���t�%��sd��̻�~E�
4�Pi�1j��~�-,�H�p=:�G^�ڈ3��6����%NU6���@ ��E�a��o��UJ�!�eE,�I��zZ&�y	����ѿۼ��U�J5��F��c߳ s��e����7+�*�>�:O��#���41�����g�βC{����^�?����8�a�
}���MF0����C:�u0�r����}ŊT�J�l;��6��|�@$���I�ݽ�w��ޜ{��km!)ƱX.[7N�1X���NIh�Z`t7�Z�Τ�3�(��l��U
2޼��aW����vٕ2OEj�!���d>�:�dI)r&��?�0���D���zE]IPd���\ ��U�x��|#
�۸�N�f6:�b��8���)�I	dEk���}��-�܋�-�W���GA�̢(c�J��z��M��U��1[�~�� �i>�ܴ?��V�܄�8i,PB|K_���ذJ�j�g�qpWC4-�Up����-١w湺�H�ةb�)#A1i��W�3ESt�K�� ��1z[Y��L�!��)�K��|�R`Ŋ�p�aU�dhùh�K'_�6�E�;������� ���y�"�_���|�9��Ik_�Ϙ-Ó��!�q-"*;�v@�+JVm���e���s�J�N�s~��P(�ah��v�OW� I1�c�h���l����w&�+(�Ƶ$Q,�K�����B��.��f�I�?���.s�-8|���K�y<�;�7˕+x�).9z���e@��@n����l�ڑ�&��<\5$o�DxF[zF;�]L�t��4��f�]5)����ek�)�0�ak���lT?���	�]
���n������H�2��G��V��)�7X���1p���6�*�2��<���r�R�G���M<(��I���f.g��{?�:u��9�_B"�=�Lq�%�u����fS6Hc��@:@�ܔ,SL�IFQ�p2�	5>�Y�9:��9��o������|�a."���/����P�����?��cyj����
ׇe�-�(��JN�~31��
���ra3��a�6*��"G+�/��H�ηT_�0J��:�����%�RfM��%��TV�C/��/@�y��%�VN:�E^��b�<��M��E�im,F�c�`�7;lP�>�U���$F�?�	K���7�W��;چ�}Y	H;���(�B�� �8yS�����L'�y+�	�,ٸ�0~�gBG���z�0�َ�B��t�G�Y��uZ�	��3V�N�6	b�s�#�o��i��;?[/��Or�w3�ű�53
�ҰCB/�{%W0 B'�@�Q(B�0��Y~�����
ߡ��MQ��9k��#Z=\r���,��5�O�b��D{�v�~؅��7�6���Wʬ�`��_���V$��Z���y�]�3���Ĕ΋��,W� P����f����wnh��=Nrt��pz7�ջX�#x�E��5�[��n���u�8J�Tmꗴ�jp���n�J҃&��,�}�q^Ѩ9�:��fԊ靚,����	ee�\�|&�Y�:�E�X�~����	ۅ�8v�� �b�x��LO�W�`�_ف�#S��ºܲ��]�0����+���C���MjR@���G�h -�Xg8�qf˩�_<yS��ϭ׸M���4�آp�(e/|c����ƍ��Ι1?uDi.�7��q�I�H�.������X��2��G\D�X�ə���l�	��i�
f�,�v��4��jG��ш:3��e��]�T�s�A�QZk&R�>?C�����ݡdM-w�%N'�W��>D�8R�M��u�#����������0���g`3T��	��1�B\�]�9v[Jg-��d'hf-�L��c̐� 
>J��%#�E�Ub�G������C��MK��E�6^W��*��)�����m2��$䩢�"=�H��ԑ�W2�q��\I4�sgTZ��<�js�8�Ϣ�4C�Y���k6'F`�e����� ��</�tԣF�z�p��l���^sޥ�A:-jH(����X���PS���_��y�;xH��ܕ�2�V� ��z���a�D�mMOk�J���c�%�c7��������˙,@��\�r��{��k��F	�͉!E�k'p����$C��^X:���V���r|?��ώ���K�X�Pc�����$; ��""5G6ҕL)�0�M5��$u��q��=3~2����S��1�N� |�G�+����{�@6_g���w�'�p����ث��IE���(H| ǽ$|���A�P�$��w��YB�VC`�o�۰��k!F$�I�vTk0�	l��処b|Ҷ��+�.ÉU@b�J��#�;b��$0��kK͘��/|��Ӕtv�;�p����[�)�\�n`�(�kF,e��;�^�f�4�Rw\������=��u�2��C /k�)P���h~�ܴ�J����h����ۛ.Z�%q�2�CH��!ƙ��Л���n�e��$�$I� �(D8�1���"��"�.���n������,wPK�K��s���C4YI��1{8�6M ��V��H�f &jj*�}��z�7�Y���J�ɘ�J4�Bfr��U�j3���_��貂�֜�4n����ܫ�	��MgJ�!l��K������e��Bn�I���R�F<L�t>ޝ�>X���w��f�|�������{���z��od��$�rW� Oz�g;"�+��|�L:u`����x���P�u!R|�]F���WѲF��ƌ�f=�Y�b���>.�V�p���ҵ� /O*�H��ɲ	0����$�?Y�,�d�[�����?�ʽ�߾T����vk:@�HѾ��R��6Gw�cvD��*�K���A�g�k�lH^�]�c�?\���_6l$�{��y�Kn�&s�l�`:�>Z>� ��q~~��cK��^/枸<j��H�$�u�Z����gC�"���i�]��y��������ޔd��XFe�!K*Q��#�`+P���BH�r�T��`�p$�
pBt��H���ah�����̭l��ƃN�Hb�W��U;xX�=H*�����N���V�%�p����F�Y1�4�{(����̀z��%�y���=I�4���gto\3����q
MP)^�w���޹,�M��b/|��nR�(�u\2�b��=�$m��̭t5��\['��醢&_��6SY���6{��}V1��4'/nґ��3��s�7�}~R���-۵�h���f��k�FK��adT���\9�y	T=�66�x�&�f��)\�ۍ.��;�گ�t�o���X���a���c9��J���@��a���jOL𞴢x��)�T)�=r����󁜧�S�(�%A����c?�"���:�����\��C��2�j�9%W�[����I� I��ɐ��:!�$��3��̱����s�n��>���+g�63p�e�S������p��Z\Ԟ�ܝ�B����1�Ty�Ǘ�n��Oy�ɾ���s�[�B�ۂ$5�x�����Ӗ`��C�c�X���|>q�X|Lz4�P�[K��>�z-����kcG������L�����/f�o,�덈�O�����[�����2�njR;�� )��A�-F�)��aUUP�_N���5Ln���̝F�{Nx�B,�z%��;�@cv�%�˂���̫�)ro�^�d}�+i���Q�Z!���{M�rh�;���x2G���z����F�p�zo^EAJj�1�"�����WCt ]\w�l���p���	��l���ւ����a�j{�6m����xiAPU��������1�wm*|���;�B���m��\[�B��8DW�
i�k/��(m��Ғ�D��ج�T0#���^UQ{��o�G���c%Y�s�mH��ہ�����l�3�{j3#W����=����Ah�0J��	�]ͅ[�-#�|H۰#�V|��}P�_��U��o$T��!Ư
bn:�.��v�MU��7�8����f��{i���Q�Mw��3�˕��=D��J[Z�"w���K�GC�����X\��M'E=�țp��~��%�Qp)��P�W�o`w��Ͻ�q`L#��� c#�`UV!ٙ�S�ު�fk0J�����Ʌ��M�.�Ac� ��.�j�����LhE�kk���٨�PǓ����!�+��U����E��"�
�
��GK�4f|�� {��0�0� |l��:.[=$��h��'&�8��ǣќ�?���a�X�^L��m�F�}� ��h����Z)܋A+��{�.�b/ߏi���$2p�1���? t*������/#	�B�w���_�-U��נ��dܩ�&���?8������mAk�s�O����w�9���H7�'e�H]��8�6FJ
�{~���h��a2��b(���a���])a/BZ��}�n�P*Ҟa�l��8���� ��*�꙾��S�\���t:z
��a]��; �[|3�pS2.�L��{k�N*^����p�q����ټ<�w\ƔD����nq-m� ��4O`����2�7��=lZ&�G*�TÏ}�w�w��ܶ��~� ���d606eͽ�i�F'w��wv0��SA� ��r�-60�s�z}s*�o�CL�����J�o���$�����B��W; �p�Ö �n���X)�0g��x�%��g�֟%3D���,�lC�tۃ�ǵ2��#�?pv����<�Q��3�=X[W��R-�z��#Q:M	S�i�̰�.��q��MoS�W_�..��j4X���H�Q�	s�֤j1��v�~�;�7��u�2&z�tqf�ԝ�k>����P�/��Ql��)��~��o+T��1Ρ�n�\�1�Vr�A9�/���>�Y��\���a`��2t�8��at�ǌ��d�e�V����}l㌣�q��+$*!5|cG!GMW�7��+�H�֭nӣ�=+{HAA����zۖL{��幣������R��T�Q��̕��v���Ȃ�P���P�bœ9$M�?/]3Ԏ�OZ�FH�����RfO�+2�2��r ��f��Ƶ��i�:4m���
۟*˥�C��l�]�}:��6G�x���_*�Ah��mq�Bh���iU܂zRm5>I��S�j!�"RS0rP�R��BJ���B��#z�2�rz�_�F�Q�S;jd�2�i��	����kq�T"
ˣ��}�@t��=����Dfc���m�wy�U:$ɚ[`�gkb�pAIw������Q�5�@�e߼����M�O�[�������^[��<>]��;2��C�](p�cJҵ�W��pK��B����'߶�L~��<[��:�<
��,<�{�F;����P�9�G����!�:�%�lDbOw��P;���8t���	K�e%���j�ss��7~�y�����<���x0;p2���)�}��qjA�&�3�HR�k!"��j�8��7J*���>
`��/�*�ea���
�.lC��㏳L�5RȪeW�� �f
}��ͬ�#�('Y�ˉ$�b������%@�U�%5ɮ<��~:g�pjI��]��}�Ԋ���L���J���H��M����+5V�b��|��	�1��T��{��A���݊"e3�Z��zH5LvGR�tPt�?�BR��?W�����I�S�
p����C蓡ojL_P�̪>��x�wа4_�,.N�@�4����!9��.���Oh�ƪ�Ű�s�~"T��r�*���I_�%K�<�L�1��:8>���>�;�@+ڶ3P�zvmWH�Ph����c,��ӉO�((�kv��l"��4��;B��&�N;�d���?��lR�xy>���f���c�b�c������6��ͻ뛶�E �MǬ���'lf��MO��2�ȼ��yMs����x�T�PP,1"*��>)V�?e����v����툏N�B*�]h+o��ޙ �:���Ԏʱʫ!��`b�ᬨr��*�Rp�Q�}����e�w�]��sJ�}���s�X��y\�X-K167�D��NӀ;��5�Z�#�wVR�8%��"���%��L��}x&�J9K�Q�l3�+P���.wb]%�Uz����B���D��M)��%�_�7X�Ӕ?�o:z��(��ȩ�� K����tKtDܦ|peH^(�L�l��a��:U�����x[R+EE�BtH�O$g���,������������OZ�����Ixc�#6��tlE�Z^Za߈��uB����+�R� ��d{x�&��'����#��hFe���wen�y��V"��������5ǽ:M�g&OD�{�{��H%�	Tp��6@(s�4cA�`  �G�����=����]��������{` :]=$�������N\�|���O(�6l�HMx��x � cذT����p,�Ӱ���+�� ܵ5rN�U��E��h�+B�e3%��v �{���bvV�]./�ԚF���MV�9}ʁ���x0U�PF2%��1��H8�=&@��4�\v����������v<��Da�u��?�.J�r/,�TbaPJi�mҵ�#�$^�2�GgE��]][���g���v�z^Ġ {�?�3Ù�ٹ��-��d���qrM�T�
I���~ԙ��@�"�v�c���̌Q���~hњucS�+|��w��sP*������7O�Pd9�;�*?J�->:�ȂsÃ���Vq���O����M:�<��nWh�s���|cV�t�epU�?��FZ��'�	�i�8'��)MA�x��Q��c�`Z��a�!G\����ӽ�;yU	Zo�Pke,^�'��,4V�e�ｚ�Z/���'Z3�zCB;�������</�l�2��.A%�����͉=塻pS��bb\�d%P+i�^r�#�v��	t�Tef�4�Ж�� �)��4>)_�R1�?���1��L��oQ�v{�����{M���ւ2!����%�\`W#<��"y���S�Pt������~��z+���"#>Un��[TCk�A��j�؊!Ȩ�
`�y=�S��x��3����j����ù�]!ge�VW1X|b]���t$��vm�9$�Bh�r3�tʾ�o��&w���u�?�PN��}p��$i�x횦,��	�+g���g��W��ݦ�a�#��/k���3+%�!�~�-~Mt{����C��ٳHD�;��R�w�'Y�g1��@T��d����,�a^2*}�.��7:{1״�s9�nz=e����ӳ����00V��%�;QZp��P�w��hr�n�bQ�p���7�Ҫ h梨͐�sk�2�R�+��aF�4f\��$%V��jt�4N�W��������EM����2��*Oy���h�>��D3����KӸ�ͩ?���ȭ��cA��~�J�\��J$��44���%�O�|�-1�0�nW��h�MfY`�z���Wc����}��=}�4�A��R���,$,j��Ag�I��Ԯ��u=��>��L,�-E9pKLZf�<M�6���oWQA(5�?�0VQ�ky��lA�`�v��Z�HE>x�m:���j9м�o�-3�Yl����`<����Op�4܁sn�\�.�R3��)�T.f+]����yfq⥺�歗BV~ʳ���2�+���V}���n�r1�Y� ����dR��	���[ 3����s(~�+c��S�@�d��Qv�M�	X �C05�l2d�N�5��| #焓��I�u�&��O�6�x�����%�sZ��
�E�b�C��஬ba��1<�{	3d�Gn�B6{�s5�AB%v?����&�@B���*>-���F `�SI�T+9����>\��*mʤ� �]ү�1��s,�{VQ/��3)Z�&�4ގI�mb��fw�G5��N�b:��f��Z4Ң��B
r�?�?��RR��w��:3l�s�x>q��������[d*W�%g��Zϰ�,�!E��P����M2���`���G�Q�[�'X"�v*t:y�� �]`r�R�h�/sQ��Ѐ{���R��I�� 2p���FT��| ��,��긴H����.��_R>W@f��+�s{ �I�rB�*jPQ�>���E��(WOk�}�d]�#��(@�^I��+����+�يe�2c�J�E�r~b�:���k���~�9��yFD6k2����K�Nϐ��Vu0l��EXf�%�X���v6��Ho���;�´�u���!-��?��I�����(l�+1������]e}c�݉ea�a$u?p�Ԙ�Md�}&��p��2nJ�<���B}���X�����w��c�fѥ�PJߦ�b[!��)�֩�%�9ٰ~I끌c�`E\�Ņ�Im>�t�D����8)5^b��+`��@v�Q�����gz�}�1Y�a����g����Nx��%z�̑I�+��<l_�_^�A|:�X)��F�e������t��Q(�@!�C�ݕ��^qO��S�T��H�%���L:�?ۀ���hE[��vO���莽;���8���ai������zu� �[�UeQ��K����۰�f�����u���2C���&�uM��h�z��v"o��s���\k���p:�.1��@��<L����;.O,� ���!���� �[~�)�����}�	�K�W��r^#���1G*�jxP�	U�!w��f!�.�_u����y��
�>�r% ��ΐ����Ygr0��:24�5<V|y�P����r+KA�k2�2}@ ����c�ݜּ'�q�@��V:���b�R:�A�6�}!��8�8�N���+�NF��OC�u﷫�F�P��Q���Ui�IJ����7�p�#L��y-�ͧ(�H�mK�E��	,��qҺS�eo��h��>�w$�{	��e�mx���_��a2���bKq��4��6V2>�_����~ta
,��+��l��z�S�*h���D̪؁��G�ξn�ٹ/��e�R�נ��ä��OFvr����v�=
���EF)՛K<ţ�fw�ĈC9�W�F���e���������Y#��?��ܰ�|vO���BJ�SS�mc,��"��������U}����ܙ۞W^��7�	7��O;�W�yg�-ƒ���!}���j���(����9��5ح���U����`���"']ˬ}�\�G*;M�� �2Eu@��[kb�#�N�}#rCoM���~���7:`�J��Q����������"׀�ժ��F��
Sʇ��Ѳ�S[��f�h"K�Ď�Dcs�;
��9�|���@*x�ۉ�����FX���ڌ�`@���� ���R	T�=�-U��Ꟊ�/�H���@���;���ʎ���֦y�a�W��&�]y;Tee£��ƪ��N�@T��P�=�->h}\`}��1���Np��@�T��f�w�_���4���ɍ���gV�E��0��RF�;:Zme@)�_
��s��D`��I�Y�蟞Yf|���7S_����XyB�Rm��W�,�a���e^	X�����O#�͓��+z>��W2�k9�K��e\��Ѐ�`��9�D�V�Uǂ�:eua�47�ڴpl*�z�=��sI�Lv����}�%,��$�J�
,�17jq_:�d��No$������8װ]��SW�����( �[3K �/v��;�����ɡ*�"�2�� 9����0:?/a�骕����t+3���Ო��K�KLH�X���g.mOs��MSL���R��$i�.�JY��d�T�R7Ņl��4(ւ��\�ɚ>4�$�� ������t�M�̵h�`X�"��m� � �V�[�>�փ�d*Y(]ݼ���$l4�3(�^;�"Mл8��1�J�B����`h�ś�Q��0s���ԙ��6�Z�x���L�j��8�&�lw3�mOyV�4is�"{����|��4�#	�V�g{�>z��5ܑ�|pJ���l��X��ޚ����a>5K���Q�i�<<�9)#0�zM���Ӯ�s^�`��Qh��Ū�$Ӭc�vG1^A��\wğ���
J���f<�%��q-�������)K�9:zbDk�"�:Ku��K�����k�<�@��Y�L��i=�&oϬ���[�'|QT j�ਿd����>1'��rD�t��x�����p�۷D%�H[���,T�Z(�/<36����T�Y�1o�F�"�w	�M}�|�N��e���0CF�'���"H�Q�u�)��Õɒ��D5�.~�C�!*��u���T�h��FÖn-%�`O�-��X�^B��h����vO^{F��p5���Dx�l��*E�F���rU�	NK�i\��N8��`u��;l�����ȳ�����(m{t�����x���T�~�M=�EƝ����8LVj���(K��k�������V���x�{fD~�#�����Nl��]�}ae��/Hr�8�ܫ~��F�������JrhQ�#���JCW°�۶XG��� ��LG)�rN^�E�����¥���k(JX�қ$Ӧ�����V��)Tk��<2�硿��LhӾ�1X/a$���\�'?��۽��-�Gmӫ��to-h�\E�����q�\�([���S��J_���DD����o�K�~A�I;���Ң�Q���0LmW�)�1،/�8y�y��.70��%fV��@e��V�c�qU,���e��PA��t�o|��͍#Qf�[��<�=e���)�_~V�DB��Y>Nni�!!�G�G�Ζ�]�"#FI���Z��tB{�d�"l
�F�+.S ���0�\vRt*��ӛY6�L�<y��|�=��!/p�gqV��p�+�v�^-�M���t��6�
ʭ��挘��^)�Zz�R6h�2%į��iwj��۩�\�f��+Ӱ����������ZT�ĴH�]�F7�,V��Z%RL6�ۖ,�i%���� $c�1X����mNe}�n���c���Z�����]J1�-"��s� J
�[I���Y�Z�f�K3I�E�&���t�g�(L�j ����M�6�_�s���l�\�?���^R* �3��=���t��J'���P���%V��xC߅R^��E>�Soյ|�R�}a��#��F�(���H�֌���(~�G�~�����;T�|͈���C �3��x j�`x:\���ȲU{��U�I����>��,��W�uu����r&@M��eI52�'��iG����y�Wt=A
b��}M
��&5E�m��X�$L<�ȣf
�_�vh�%}eg�$[�����8>�3��d�W�8��l�*$�/_�� �r_��=����^5vH��hV�5\70`�9⨦^��c�E�h�!�hn��4��r`fz�<�1��S���N�/�$��{�jV<r���H���^�ޑC��>a���0�G�
� ��!�ZP.����IK �Hp/� c���$���{�BB����s%Y"8Ԧڶ#���q:��}��]�g�����SSK/�ys�z�W�*d"p�^��\��-���l���_���P�������V��Ee>��),�&.'�\�,T�S�Y �H�#p��et/h�hP��jI� ����Js����M���ڇ*
՟��ݶ�4V5~T��X?]��K��:�uP~ OR�~K��0�u�3�^�*/l�kC� Y}�5���ZFN�D�K��F�>�k��m�'��a���`2 �JE��890H�'���B�3:C�����؞!L�Cp��\K���ޥ%�����?'F^�����G~=�T���	�;Q5�ɒ_�sD������;9�[�~�b�%ԭ�ݲ��,��pQ����R0���V�-a�9~�K� �	tk�2��6�-���7B�?���Gr��C[�+C�=.$l>�lܐn$:gI���\(��2�E�ݓ�8Fxӵ��oRKPD���ᐩ��14��b����t�`̿`g�]?� &�7��γ-"ղF�v��+�i��/E9q`IU�e�呼��̽�,|�����X�<&���p�-[~�AE|7[ ;�(㶦�	�&v���Q;� E隸�md��6=)(H��T���'i�����s\��u�]j|6W��٦��U�;!�i��{<�����蠴ڜc��|�3G�0��U#m�O�����Ex�1Se�;U������g����� $�:R�[��i@0�<S3D0B�:l��鲩��K�#���n4�Z��,R`��̓+����v��v�KGg���2ђ�i�� �w��s��Μ>����m����G�V'��q���7׀;�In~�{�:>�0r�5���8����iF�#~�-0v,��iJD���M�Oj�y�ti$D��"���O<�� YL������F�v^蜙�d�e	����<dzH���S����goG�F9�)���w���!Q�'��^�w��Tź��c#�3�eQ���D�~�IcՓ4ML@]=/uӓ ��N`��3"����ԖR�?p�m>�C@p1��M]�rg�ŷ�Y��wZ����4���FO���S��q����qg�[�Z�i��&��L����J���Uh�ܴ�&\I�D�� ��\,��Vb�U�����o({|�����ΡϨ���k�&nhk6�V�"�79_:���9��B8�Ⱦ�݌'�Gh*�{�`�H�2c*��͎��2xIL�5�R0��_�A��TF����j�q��~L�~���h�W��âd;�*&Wjp����mxL]���`�Ф|~��c�H��e��p̑�Z@#Rۣ�jw����=��0r\0R⹢m�"0�\K��+.~[�SA+��,)��y�e&V��ݎ;����,�:���1����@�*�!�>����j���b��$�_zX�r]?n�ݧ&>�T�-{�I��?�����Po�˫]�Ą��x��!�����`�Q����]Q5.5�L��,�ReU_��1�_.�͑����=-�  ��~�����!�t 4��P��ew�)�+��6�CV.��#��4�x|���ˇŷ�^������t���3����L���6��5�jP�:m.o��Xj���|Dt���}͇�Q;re߃cA���ʕÒDMM	jh�k31]q�-2��<�A3N�x��j��p3�İ%r8��Fշ�o:Q�����\�&����=dC��
Fcv�O��^��ÏY�ߙҌmLL�$%يߞX@D���'��ə��� ����������(L_����i��Q�m-����6��[(���U+Mz��R|h0��6�F�۝��L���Ԡ���=��J�)=K8�"�25��������`Ԫ74��ԯ[݋W�����n�]�.LT	<E�uL�jp�!�f'N��h	"��o)��_���K�끐!�ыw�Zu��B�.M�"���S��G6[��P��{Y����ڟ�->XYF1~Q �knB�}�!s:�']�|���ࡏ��n�H���I���/d��ŗ�]AL-��&0͐�����a=�㾠7(���z���r[�W8����j4D�꘠���y�D��Ѓ�ܨ��%b!C���M)1O:���r�Ǵ��^ꍫ,����;��o�|����q쁭׻Eko�
���ۅ�ٖ�3 ���݅6�G��;�G��K^�v-*6Y]qC��k�˄�d� J�#��f���D�����\�VD��K��:�c�,�΂��&�W�~��C�_����wK!]Y*4 z)�5bT�|�2$T3��_p0q6oҤ��2g.�D�"��]��>&ޢ
�iJ�G�K߇Ҙ|���%d�1e���VQ�;Ma*$���6�5�3��sC���Gͫ��¢��\�^E�Ƒ26���ؕ��H��,��ڣ����Lmֵ3�"��i:�o�ݲcT�́�:ϺU�mX�q����v��|�'�-�-MY��Q�Az�w�p�
)�n���m�k�O5P�-��Y%c���%���k$��H��ww���p��%y|&ц/%r�s.��#ZuG�n�#a��J|�w���=�X-�!;���)	����]Pj�MTtI�0�ʋ�v5�QI�_0�G�;/ِ�F�1!5�)m��|)�(e,\A����nw��/P=l��ݬ���[4bU������ �wi��<���zW#�Fz�?�A������nf�}��!+��4}`���UQ�=b��1�O�X��6�&� �s==�e p%N�m��RãBb�mF��9�i���$����{�S�܆6G�d����Pm��Oc*b����|}x9��n+�r`�d��Z��姸�#xB-F!�����܅0�Iڭ�߄J$
�j��e�̅�Z|D� h@}������������e��a�#��G7�p4���mg���K@�Οݘ?�|����{I�I�ۅ!Q� Ω���[��>2�&T*Oռy^��|C0,��
1;&4���� �8��p.wo�:,A֬P�����k=�.d;�dj2iLľ�Qڵߙ'�=�5��a%���a�B�:�B��f#�12�<R�����8�y�JEi�*����W:a?t75�Z���L���R�,���2�d�(j/�
����>��I�V�wHw�3*�:��p��x࢚�c&@��5]%d&�ګ�V_�Gu'�G���)^�b����F��+'�"��m�؃��w��N欃D�N9E�3��Q�N�<��c�4Y�p�gվ>п�+�ƌSݾ����2�gkZ;ƫA?o��۪A�������'�p7�k*�HiHRA=H�zDk�2m5��zm/s�6�Ӛ�!FU��*UuW ���B�i(+?����kɝV�)�}ƙ�����B�v��Bܦ\��J����@z��E=�~G�����
�*E��!:Լ��mh�ߗ�ֆ�缘�m��:Rj��\X��V��������̖�:cD�0��f7�Ɛw�o�-+�&ڂ"�78{��B�_��Hګ��o��@|}��ʏsuE���3p~��~.`�K*&��#�W�Ζ�ٯ33��/�2�P#n,�'\�f	��jSF��ӥ���r��ڣ�k��j�L��s�F�Z�4S'o��z�[r`��4;��_7�"rp
��=I�zƐ�i�qң$�)��A\cD����"چ׋	Wĳ~Y��ˌ�hE�;�V�5<���x�3���7�~�su�S���Q�5F�H� ���׽$���1��g1�I�aQ4���26IJ�m�QH�@׳�8Oz��Mz��A����#O5���T�α-���A��m�:
Ŏ��P�Y�]���oȺ~��6���)&�_�(���DS�[:�`����A���˿�9ӿJ64��7���U$\)`Zq;{4��t�5��9�9�k�� ׸��s�zp���"̆�{��ӛ�$K�d�V�_�f�U�QC�([Nbg�qDġ��uXҴ������1�ݸ�]-���!w���q�<U�ʀt�	��I̠p� 7$:K)����+��bo�ԑ}��8�m��W��Wg�� �_K\9aP��>���Ʉ��x��@�Ib'�$;4ڍ�E�K��xq��&��#/�R���D"�]�q-:_�I���f�]��S�$[մ���)ۗX���)�ld�^�Q�����G74b�[�4ar��|F��
���}�'с�-g�j��o��93u�"�����/t�����~ҋ㬪Q��x��>���i(���r(�%ҟ�3wW���2�8MFFupf�,�t1����k�`���M*���^�L�b���JU{φ�u.���U���,��_��C$�Pr�E��ѱ}{��/�y�h��� �^\8�t*��1� vLn�Rh�"&��f);J� ��A�w�o��6eQ�S�]�,�Ӂ>R�F�*g׷�_�-�
PŁ�*e�������1"��hR�`8`~ �!�t������㽙���h�} ��u�&�����Q.�p����;�{�:�
ġ����e��\����'�h�A��Pl�LH���C�����8��ݵ�E<�n���wr�`�H8�4�JŖ��!�s$.۶t��bGG4V<���%���������1�ׅ����A!�>ts -�l�b�n������Y�̍��Ww�|i?L^��Tx���Th|�� n*�X��e-��(�� j��S����¬R#��E�����K�@Π�)\Gi/KJ�e�ާK\���t�3;jg~���,����#�>`��!�ò�Y.t���x����I0������S�~��$9��;��C:ꛝÆu�ȵ�h����ks	��%�4g��c��d��0�Fx����\�+N_��o���M�Y������$Gij�b��o<�儹�uAL!�E�nEʯcxu�P���\y�-�-��Ӎx��_r�.l!1�ށ5ՅI�z��J����Y-U8@8����sf�j4g�ǧ�_S9����W9���j�%A<�Ԉ��RBZ�'�+H,
�L���o�����X�+߇t�����f�T����)�p��C��GuR����h���B�����~�P�}�_#�֐�C�nF#�W��� �g/O�f�fFf�������S)�aS|^7[Y;��������J���Jx2�r��*���C̙���ݜ�J2�ad=�=���/q�0@M0�.��WK��͙Ŕ�X�:=Z�M���5|8�ȯ�Ť��Ks� �Ѱr�Y?���jӍD@�9�7ا�Z \� �8�E���/ڵ¹w�ܷ�z,qgtˍ�P�%�C\��������^m��t6�B�	~1�iǪ/���@_��*|[*t�=��*����G�a!���&�[�]*��M�S��ޥ�萕��}���G:%�[R�UIJ�����e�kw9+H°S��o���v�^'m��Fwz�M{��k�lv"B1.�O���e��f���Z�#�	���mt"�W��������8�����-��$ED
7�UƄOv!8u�f�`4���d��K�\�;
H�g���5n�6`��U���l~�W괍�X6��::}��/ʇ6U���tk�J?pGƪ!)Q�����qͻ��gb�o�hVG���#s�ܚT�����cܐ�Q[����OgVj�D��7MבM����"���~�BD��=�f~�/���K�Ԇ$���:%ew�#�ɏs�#�j.�����Bz�/~��;�0�?��QU���|4]>�����FCY������]���5�i��f���ُVG�9�_ŕ~�W�V��X-t�6]ė���8C�~���|"�&�T���CU�x��]\.Ie��@8$��hhe�i�����}���)d�ӹ��Έ���X���=��avW��\sC`ϳ(>[r�D�1��Ҭf����h\\�0_���tBcӶT7p�}��vf�:C��ǰ���c� �����G���Bzou���{eo��T�6KH�BfTY��~�*��pG .�ϻM����]�%�qe�2 ��ۺ��>B;�`�����?3��R�ݵ�s@�&��b�e���1-�O��D,A%5ɸ%p���_�'���jY���i</�,Q��Z�W��^+��X��a:y��$	�&�����gC�P�8�/k�ާ�-dHo��YLy���%k;q�蓏�s�7Cx�]�
{�`lĭֶ�'�̊�?���ş�0�G1=>�=z<��$�Si��^�7���a�S"�5�� ��A	��������nw�7Ｓ�U���)���JoS:
$�ˢ�B�h��Nܸ]�&^�M�5X��E��cZ+���xD�.�w-7� q�m�)� ;Zc�_Zj�3��=Q���Sj��%wV�$�]�����~���y��aM]�H��Զ��Pz�f�`���pM�Q�҂[@�,4�*��翊SE$�:�.����x��`��dB���+�n����#��o�h����Z#������13�K漾�������ǿ���d�D������* T��@����@5�RUl�ny�c	*�:x\3���}&��"��{��q�FK
�C"~1�Pb�sY Og�����,���6p��~s�0��x�"V�_��9����<�@��Z���K4�Vp�
y&�ر:��v��Jܣ{�����gub�[aչU���
�LЙ�jt��� Q�Bڋ�,S5���a�ڿ�|b������2��H'��}kz�</��bn o+y{��ԛ�6����/���R͈@����ZթH����e1@��R��&j��G�@�&�ջ�� 1$��փ�4� 6��;V&����7*�DH����G���\�iW؂����|M$QA�[MF�'j���G �=w�|!I����!��A߲�a����Eᴪ��k8���fBa�C�MZ��
�����
��q+�dng�#� �)M�Lw���B\LR`�7V|��y�2:�`�V��$^�t�����֬�F}���/Bݯ�Z]_�����+ָ�ۯ�+�hd	i��!��V�Ú����
���7B�v�o�ѧ��8�pNC������ Ѣ��j�ǙT�}~�B��}l9<m	���" ������au�Ł�K�:�4����o�9
���//�B���	\��,�^�3; A�o޻�o~$4��������G*��!��uk>}?P�^K�v~�&E1���-��t�����$36v�����&��_�ⅎv�t��e���wb��R]R2���W�o��̴��'���bT[\z�����,"��q_���<%���Т��ܠ����%�������3/s��a��~y�Ql�d#����M$���?�rq�D}A6:��XlB��j��,R�=mzj�P�Ϙ���Vyx`��N7�O�zCu4혜*�rO�]ј���ɥ����P\�ߍ�s$���rB�5K)[��=&�����к׿x���	�����R�j���U_��L����`��D��%�"=���Z�$�m��pN�����	g��i�3��%����#��P=�QH-[��+��
F�!��(����z�?�,P���I�C��d��f��#�$�}�Cȉ�[>r��t`)�M���|�$V��?ȧ�FX�<4A��.�cj��9@w����sqZ`�"�=��/���m_�1�b��?��n��g4�%b�)>�W�a$h�������\����*[��.|@�/�"�W9ĸIɝ( �!h���ptDev5�^��)@͛�������@h$v�դ�/�D_W�o&C֌!��SdO�Jۥ4���Ӧ��j�ao�i0ǋ_�����)]Y�<C��̓�����n��B�MzU�N39�i�� �қ%������F<5��w� ���@!�
����=d<��@ ?��8��Ǖ��AߧU@CO+��:36��K�To�\���DD��q�#����7T��4�;�?Q��v��r��)�χ`�C��x'8��Y��{��Ԡ<�E~s�"��3�c�f�.��Ъ��2���P��OĦ�4�/�|��������L��@�Ε?�$59��d�k��g���m��
�9{�1��*$/�U�UNJ���d�B�&��Pbq��N?��x���>͆nt�c�jrD�Eq=i�>i)f���G(�j��`�5M�P{����Ӵ�1jgĘ�%���D�<�k�'{������?��7�7p�/"yjފ��U;L\o�� �.g�@�)c�3A�����p:� 򕁫r���%l{~#�}d�����r��ͤ/{���;ڮ>�L)�-"K�4�zҁ;.�_��4�_�s�B�c��B0��U��Q�kD ����L���4˨5xL5a�t���Z����_�hP#�p��P�~�s�S8L�z�A���u��-��8zy��hy�Nm;�m�Tǜ��������F���㏅��|���p������^iߔ�t���\aB�ऱ������C�+˄��m���n`�rv�ȿp`�tI�R�� 5%���
Y�5^W��݈��+Ӷt�ĭJ��gЌ,�~%%萝OI��I(6��8=q/�S.��*�F��RkP^5,~-�`4K�_��4��p�:bRu���o����M��j4�0�f猒N���w��LA�K�1xF�h�$~��wj8éX�S=i]�a
�X�⛐�əxv�L�qH]����z���.��Ok�>�bT���f�D0ʄ�Վv��`V;�l��w/:Ba=��(�����GZA����̜�Cg4ب���9T��[�9�'T����y�i�y5��WÎ�t%8�eu[�o��m�ֶ"]l��}�{޼	��=�v�)�Fa��*�6�T��f�Z��VF�m�g$z�����n�h�1�\�h�c�a�*���C:��I���!�XI=�3^��W���s�X�9:���e���:�+f\{�Y�5�~g }'/��bN���E�`��6p����Q�^pJ�c�YTn��O��.�,X����D*ѻ2%����׈�&ܡ�2�9��g��/��iӅ�K��sc߇�]��HVl�6�=%��l�,�H&-U�kLM��An���z�����1ָZ�:Jz�N�G�-��|���3���[Ȯ�8>휻��p�h�r:�r����}���R����4�߂I��3D�+G��W��e~9'U* -�>r��Ł]��0�V��q(���H�":c�.��5�q�BQ��ۢ�^\�ω���>���9�E����ױ��h�Ԟ��M��Jya�Y�����Z�٤���;�7Dd�����l��b��^@��ï�eϠ��f`!���O6�+'m�3K�bM��`9Ѧ���Z�N��d�� ������Ax��<"�t�]�K�]���� \n�A���\v��86�RJ<p������M�
�w����8E��t�(����r�J�W���8u��>��v��%Á�P޼��ɣb9��M[ǥc���~�<����~?!���7U,��BI��״����$�e��ް�XM�֞}LH1"�b���`��~��ӑ ��>}�P�(w�]�g!Vt_������RB���|����hC�뜮�4+����&���p�Nd6�V�ɁKO��9y,?�90����l�ʝ�68̩��I��n��s�ףf����|�趧�!�+ܓ)A/{�s��ȑˉ?��P)�4,�;:4�n���)��eW��H��\pi��h��K�����?+�`� ���dXR&�i�V�O�aay�_7�L)�S�*0�K2�JMu3���
u��O�p��zy������� 's� 3�Y�����!6:�!µN�wc�d�|�Z��C���B�T��ʔW�;O�~�/<?$����]0�'}ש1aU��fח��n!�����H��e�ocx����'��Īt�!�[�qT`0�2,ehM�"׭����cN�h��<�\:M�'�O���-����_]EQ�R=�y�e��e�9���C-����/�B3o�j�!��	ʘJq��L��Δj�����]re#G	G�A�f���;�C�O�P�0���9�A��`�a�=��P�31X������͘L�Ss�(�n�-�${�/�6z����`r)�Nj,�-(z�{������C J>�{륬�%����)�&�"��|���gcaΙ��a	�)����^1B�T^X	 m�I3�h*�ʛ�i!ZM��>^uY�+���Yd��\�ղ��������&/�\�E#*G���ŕE!.B���X���W+�m̯|��#�^J�����N؏��P���.������\;)�d���R���<2�^����.��MƐ���%:�.w��dFjny&No7���1��~;N�g�3�g��#���l����fß�@�'�Q��>��e��'ꥇ��.奧��''�����B���=�� 6�mC�v���Ts"�y�z��^Gej��jᶾ�*�Hߓ��#��UF����It�2X�#����$X�XA'ʖ�{lL).���!{��9�wNĀ,�Ժ����z����֤¼<�����퓅�p�ߋ���g�Z� ��;�>��uH��{I�&*-f�J���-���Ǧ�ݷ���y�/�j��d��l��oJ��UJ�9��)�%SZ>^H��M�)@�W��/���!��K��L�g[<U�S���8.��];6��A��f��+Ff�����|����*{��ڪ�ߧ�,���Tдw�WI$�A�����)����|I\	�X �x�����B�}�ȹ�U���Kbř�K�p���R��&�6� �0����׮N�~]]�-�p}�1�8�nd1�Y )�[7�QH��EoV�|]\\��1s*�%ej��Ǡ���m��#S�$���;�8ܑ�!T=f"�wO^��á�ή�&!}P��<GB�$���yi��̫;��W���Z`����%Q�!�?T��}��b<}H�����&(%ضO��0�=b�qE!SV���A*�/����%�UYI�䦿I�Ůx��#���W�@�~g�ށ;����qV��Ϗ�L�*������?��Q��fwE ����H&0z�z���z���b�D���*1�D��bK;�>'W�4XƓ��Ђw��cW��Ft~N�����K��e��腛&j�5's���B��}}p	��>ppM2�֯�7��A�}�R4c��|���O�  e���}��W��Tv6k�h3L�����~�}|=y73���E#荤ڷ�k'g-��T����g��IF��7�Z6*Ѽ7���T�B-��mC^t��7e�QպF��jJ̐� �9caX���(���ܙ�9ҥ�ȃ���.}���X;��5K�� �����|��o;��	��V���H�~{]���z�����}}�;I,bV'�N�"�|�6B�q��>_�qMޑw� 5���Ȝ��V�����Q�A��4�5f-r�����[��cPC�\�͌5B*Brv(��_f�1��Ⱥ
{�����:�f�Ns�$�.���*Bd�h%��$��ES�׻�d)�l�]�}��B��t|��(�jˆ�����v�9~���NH�q/J@Of�[f�&Γ��e�Q�xRO���>�.����s���qF��o�uNq/A�N�6��fL6 վHY���������?�tҨ��v��u3]tC�����=�v��A5rÊ�l/L�?�h�K�%q�>z�r�_��=n��\���aW�!�T�H�:e�A_�j?��L���n� *�4))�T��.���in�:gu�u�U�
�]�_�[��8ZTzl|+��9Ԅ���EyQj79�E�8�AI�7/�%�c�^��*�8T~���V�4�٨�^��_��" ��`@�W���^i��ӏ'�i1�qz�4��f�Tz����x	J�j|6�ԧ��W�[�nO!%-Vzu�(hI@8����as%Do�[ϖ��Oo+�V��������Z�	Ʀճ,�ЍKL���i2B���*�ms�+�&D�N�����C4�����e
~�T+hjE���o�m�up�N�Y�F"�ӸIC�kr����J