��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V����hN=��a���)�硹<H��׮��`̼��D�g�;�mR�#rj��S��k@'�q�/�ha��pc�R�(��g�F�ו�����`d%D��G�qK�DW�+X���iv�O�O����9�t�0���`�<�F�2MGJ�g_Ю3����Na/��4-^}��ru1������>�9��& c�dN���(�lE#���f��;�B�+hTy p���E��<aZ���m����t
�_�F�v��f�H�R�5�W����@������c%���ɵ� �*R�^��%�"�µ���&�;�(~aR���t�|'�̀�Z}غ��]�V�֫5�ڤ)Vrյ�O	rR+�q�������x�7��r����5[W�k�\Nr�ы��W�[L_�h�Ж��I����g8�ʪ�9���Z��2�;1�k�:���.�j�� Kꎌ'j��ZN�u���������*�[�c8hG�	��G_���&f��Su�N�b���DQ��Z�r��|/O�w9&�[�BY�EW��ѽ�i�o�Z$w�����(t��o��]�Y+U�L�P��f��Q�ٽ��w� �e� %��ӻRp�f�xz��4���˚�2��(K@6���8e?'��U��OדGL����LZqA�\_��촌���G?]���uL�_*��~*ػƁ6�lb}���Ӟ�gz|����͔�&���W��A��O��z2<;�w?�J������2dm]���� =#K�񩝤�0ȧ}s������ ����$�a���04B��ɂhq�.j��j�����_#�"���F�X��o7P4���'�l�W��dbQ\U}����)��O��>�P�f�8k���b{��Q�=���q+�0�EU�)�o){�_����FG8�v��@;�����`��a��Ҩc�����決s�Uu����8������"�b�ԭQ�5��tnHi�%�tɅ�t���j�=���#�z0��I�mտ��>�{A��5`���B����殳 �s��(ՕY�x_X;�V
}:I�Nd2��bwvW����NUf�T�x�4����%�@΂M��?KW ��-ߓ�4� N$��1q䃔�=v�-|�d�@�b�ؘ��nPYh:U�!���N�"x�aa��8�*�i�Ex��8��ra����ɗY��Kz����Y��i�}��R�ˋ��r|��Vg	f��6|z2�2����)�e�W-V+��{��+�� �� ����KG�CQ�Ɖ��-ۏ[���2c/�����s�z%�I���kyFM3���${�������$���b�|�͸Hx��+��>�-�/L=f3�Y����q���ēD��J������~��o]rӤа�X��(�3�	<I�"�)7<�M�w����U���Ia��ǗI���%h��i�i���݋��9L����p�@��Wղ؀bT{�
g��BI����::��z!�ͤD"�X�p��*��sq(~F���[wϧ���	�E��/��0:n~p<@�2Q�f�K/ˎ��)�5TХ��سD��bg�/�o� 6�,W�k�ʊ�Ƶ�z_��w9���s����%zWe�{�($h�wĐ�.� �熦�uiS�߬X.��VeL��x�R��qkiF���4����Q�m�P1�U[ ��ymk��k�)�z�P�^ˊNd�~�ntbE��;0��6��F�X��V�Aֿ���@�j��R�ǭ��f�"�x˄=�&��:�q�����@T�hɅ�p7T3���)��J>�XO5K$�^����u�c&H���g��~>�_��6��o;]/:j���.1�#��2�- �� DBa�@�y��6YTL��W�ێ��W�Ωa�v�v����[�6;�t�%����9�����|�R��<��ߕ��Е\���L?Q� .�tx^��4��WH-�c�fr�G�� �a/���kX����e��Y-�{�}��M$`��m��du�rL.���l5lgc��$���"#�������4�.@q�_Pư=���+;_��}��j��ɦ�|�6.�'���&0�2 G���� 94>�vo�G�{ ]e�j��D�'3텟�,v�>Z�P=\�uw�[i@�c�I�b���a �������T��uBz�{D�f�5��ń�o�D�7s���W���%�ʪ�{���m>��&�b.褈���[mY$c���gm��˗߸�sQ���2���Jy�b����t�7$%��j?�^��Kԇ�0#��JHZ��i,��p��t,�� ���.��ׁ�vq�%H7�����%���k��Vj��,�6�x!�
��c�a�|�	nU8�(yk�f�)hR!��*�*��/�|Ϲ�5�˘�2�����hC6w+���ŅPx�:&���V���`�;l�E����N�m�d��3���{0�~����֩ ���O���p��%� Z0B�z��h0v���޴�m��|a��� 3�\�_��JHn�Y��o�nf��m��o��Ԗ<o�$��PNp0�4�}�"_��S���0��2Apk[wH^��	���:�Q���G΅)Ҷy���C�������{�v�Έ������R�����aqxg�����uc�}--wہzDw�bO�W]�5F�9��%uqe.�l��r�p�7�9��y"�L�~�����E`_ ��4�u^��7G"i4��-��$��k�*���b]�ED/Q��U��C��
	T�2���a�߻�����^c�޸�$"�Pf�x��ü�Ǧ(]��J��Z0xզ��LiXBZP�d D@I�ۿ�vN,H��ͦ9��e�\����8x����z�
^�=3�u�0�;��M�6x���hUu��5jT���s�^!c�`=O�#dm�t�q��a����s���Mb;l��
 d��B��&綼���Du�J<������]�v��N"�\� vU�9P\-T���}&R�5�3B|��8�����A^6�*�Q������!V��,i�O�9*F���}�+�if;LlE��R�Ӵ�x��F;��xS����4�<@��0�����h��D�>����c�շM�j)F�y/��� %��rA�?w���F�93	��f���gPo���0�
Ϟ��hW<V���<��{���u�Dd�r͇���\����?n_<0P�.��戴��ڵ�7�*��U��:q��Xk�����#��-A�"'��[��EHf1q:T�7⊲v	:�c�4w��c�W!ljҾ���<8���E�UZ?R�{��?$��V�����s-} ��C��OO�͚��6\P�|�OK4J��L�{
e0s�33r��d���^��$8�p��?�@vl�Bm������������:�v�dN�}�>q��xé���B�Ѧ� V��xg�3��OC���DZs�z�=��׮=�Q:�Y��b�e��*��*X�!xz'L��*TR��ڪ*~i�)�K�i�*q���p��I��}I�x�� <zr�% �?�A�����l��=5F�V+��7�(FУ��\