��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V�� ��9��[#��`�Ռ��j�!<�3'an��e���D�ėl�c�Exdk!ʾ<���
��rM���������|%��aC�cJl��7f��������=�s
��i��"'=�cN����"��`et�ۮX���A�����l̹�yR��l�Y%��^��QG?R��a��c�p��m�WPVɦI�������U�,z��p� �ի6�ج!��u	��k4�^�^�&�)�Ѥ�&��~t�&L��Epq��j����)=j�j��=3ʴ��!�x6�
�>'�N�����T��Q[`�v�x�	Q�݅YY�D�4Q^��/����gӇl�#�N�Z^Ԉ����\�D���?s���W
X4Jx�"A�	-a�=��t��*�m,)�j���@��ѱ�� �bx��!�b�h$�v�7�\�.�B`�M=�~�x�גZ�v �˷�!ay�%=�*�젱�����:�q����Ꞽ��{�[?�}�y�ߦ����;�fYծr�x��BQ��G`�滚{SQ1Y�H�b�ֻ�F�̉L+h� ��ʒɇ���h�f����T/������C�wpm�\RKm������e�� �����J����<�b��m�٠Bhf�?���pi��Z���`:���yg疡RS24�ϥ��E��Ŧ�N�~pta32�c(o%̧xhL�A��[�ھ���1mi��aW��W�a��o{���c�l=C�&�u���{�T2s\T/�g��y||�_�o?�?1<�,T�x�w����=�]�̈RD	��{��Мl	Z�/��)+n�{ �|H8���/Ic��NQu�P�C]"�Q�+�=sd=7+�	E�J۹�����I>��c��{�4��껄�,�tF� ɾ��t�m ��2~PhvU�p��Y�,/ݢ�x����4�ߎ�+���2� ��&B�By�qV4�X�����i�rQ��c��6�lk�.|
`LXp��<�^o:�񒒢ߏ�,J֝�N�*TR����p�iX���{�K�"�1E�9��X����tp���\�&K����ulB��G!��Ѫ�|��K!��ۡ��+|\��;���y'�rSFA���@Nw{���̴�x��Kz���-uIQL?��8E�^C���	,�c�#-;a���'#?_/��߲&�x+C�R�c'@�oj��R̂���C�N/<�j�3���ӄ�mr���bt
�ir�A��A��UC`}��%��|���%B}�8���Y�w/�ڟ:U3)��u3
Qi�n�M9�d�Grg�K���;#F�o����H,s�f�p=
��/o쪞��f i�L	}6��w#8u�����a1�]sg�o?z4��{�q!��|}Vy`��b��nx��,��i�Kp�C�6�P�n��ȣ88��icb�RA�����QJ�yv�g�/w+m,86��˓Ә�����롢3"�ORmNd��3���:���z��6��Ϝ�m5Hd�_$�3m�����߽����ޅf�JT�( 1L{��~��㐵�O7�$�#!@I��w{��#2�\����-�9M��qh���j�����z���ۜa�h��d�4$h%:�t���6�1URV��zC��OB�{��7��}�Zr#��,��mJ��8"�~�y��u'FWf�*�:=&��ٟ�9OSS��R8o�� )�Bc���.#���YU����j~���)�����[.Ls.��N�#��]�=������"n,��r�f�TË[y�LuR�&��x�ocY�ZS!e�M ��"n�g}�B�+�_$�!�����I��9\t"��p�PY��r��z٢;�%0jZ�C�����a������Ө=�Tz�b�Z�q���Y���U�W�{��w��ihiĦL��,8K�:I#o{���h;��.�#D�a�Η���Mɶ��׎�����͖ΞgЇCT��}O�&�_|���筴�SG�Cgu㿂�+j �TS��ZU���z�4p�D�O�3��*��[I�æ�7N���K��E�ꊇ��B]s�tSS_/N�s�3N�����蒀�];�͛y���m�HQz0D��7s1�ݕ�`Dv���U��]��T�H�#d�$G������nh ;�N�� 