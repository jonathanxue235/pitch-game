��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V����hN=��a���)�硹<H��׮��`̼��D�g�;�mR�#rj��S��k@'�q�/�ha��pc�R�(��g�F�ו�����`d%D��G�qK�DW�+X���iv�O�O����9�t�0���`�<�F�2MGJ�g_Ю3����Na/��4-^}��ru1������>�9��& c�dN���(�lE#s �.�g�A�|�fǼ�
��S�b+x���5tT���t��:x�'�Ԟү9�Y�A��;2V�c�8oǅ{v��Ko���&@-���V��$nh���:QM�	0�������j�����0�{=0IT��[���=��K�K��m����~l7�3�Y�5��7H$n��������q�<H�廏��-.V�.��6>�����\�������mt�4��L�cl�*x�f3ʊ��_�+����6�h��<lc��tc�Qh� tS>����X$��N/��(�#�w�=��Lt�g"��v��ɟ�j����X�������&� G)���%�e�A^y4|�k���X�T	�P)·�U�������j�/��:�;ܐf���55g�P�D>�$��?zLAy��}�hT�?���H@��L��3(N�c2X���nA14c2l7��-]!El���3d��R��6`WO\ꟷ��N�]��l6^���2�$�=�Y�������T�%��ք!��<�1�@�Y?+i��"=�X<�vƋu��C��@�D3��sj_�����f�̔�ufP�Is �$�?�|Kp����DiMh����E+��gE��E��q5e\���3�e�EfX�,O�i̙LX^�҉ �LE��YLgT�����E� �A���p�R��_��So�Uo�੐aαdl����@�7e밚ZԘ(�#1^gr՝���v�0<��=��4<�.�L�
�Q��I���=X����C�I�8���J��{��ĕ� 񵯦���l5Y �ڥ\��`.Eur��$��d�n���gFt�/�6�3ѨR|r�䔬{�!s��uh��&��n�����|`�@h]��Hp��`�Ɋ��$���I��LQ~�QU�uV1x���v�m�aj/?��	t�a,bx�ߚ�w����:��qf0���nc�8eHO��ގ^BL��!3˴�T,��F����ɣ��}�v���<DL�#��{i�ϝ�o�ٗY�r����k
�����O	:bf��a�zEآ Pݫw���0h5O��Яe=���3��p8~�rP��$�� ����&��Ɍ����v�U�L��)�G(��8��!9��5i��*���:�U;��r&D���	���s�·;Z���D��h�ɒ
�s���3c��2��i_!H�d�HE��Ǿ=6k�E�C�g"���|�^� I"��l��w�#��ݎ_S4�ZaH|�,E�N]���dqN��� f��\��z����I	}�wLg��%Ѱ��	T��Ӈ�Mt�dU�Q���"3���V��G��?�����l7��6ʩE�2�rhE��7���;�x{Q@�� ��k����7����/,}�A1��Rb�'��'���.��|��}�u��jc �$��bH5/��T%~uQ��}V�	�p���g��5�JL�Q�q9�=�-X;��i~��������i�Aע�כ{���iv��]�'N��E����F��)ݿ��S�iU8^�I= n�"qct|
��H����.�y�k׈���0>� �����ē��,�s�40h^��݉����2ίt�Q�Ͻ��T9zN<��caL��'�c[o"=�����L�̷�����dգl�"��P���(GC�7�%��O��8l��0L��W������ ˿�T���Y���w�� ��Wر����o��	L&�j���ah%��{��#2)r�RRH$��2����4~p����hu�.v�0�7��_cmFy�Jz
��&����~Ӿ�+#� ;�c�m����YR����9���|�̤��/9�b`s�MTYX�O$����u�%`�"w=�t���Q��=����L�5\�)t`KW`��ӅC�]�/�Z�@�-�:~_��p5���ZѴ�7�{J�l�v�ѷ~���KW�<��;e�.�ׁ����޳���T�/��R�#'{���?��!�P��6���\VF���Z��K �{�ӈYƮ�t"���מ5}te�O�Sɰ��u�L�G�oĀ
�~����k�%��W�e���z�sn2UVk���h>�_���fR������9(+)���n(ԲD�ȣhb5�zNq(J�R�n�o\M�@^Z[d�B��y��Eą��0'Z�8�x�x�NPl��J���p�1����	����<�Y�Hwz&�\�o���-1?�ݢ9	�9'��5D���!�φn{	�N�z�A�l	#�8�y��62�(<�b�D
t����H4�诚�,^��V�ä�C�
r�k=,W�J�sE�-�|��8G�/<��7{?�~/�����g���s�|y�Su;�k���R��F,���A��>��[h�}������_l���A���~E$�b�c�vC�T�v�������s6�*�T��)���E{���
�e����g:�	�x�c����Z��?���Ւ_��&T(s}�B�� �Ӭa����T}.E�r�l�&����0B�f�
�`m�֤��e@��d�n&�����a�E�?7��Q���ʼ�eS�_|gmXT/�HTy�ep"�v�I��QYt �a���`%�$ޖ��aׯv��\8�y�7��E" G�d��Ĳ�4�m��3[�8��"�EdVN�v@��pD�����k�'��la�ޥ��7�����^���1%�/U�J)������J-67�Q��N�Vԫ�p�V	F
��E�����ݩ��iq��<�h��%�֭�f� ���'����;��,�J��~3�c�ź�T��9����I�ə�#B2�[6�S��!�Mr�U)��&��L��������8��}-R���N\��#ݹG�R��zUT
n@�[��3hF�؉��K0��Z�gRǲ\YM��k�`k�z�_F���&�C����b!M���2R�X�|�������q���d�㱙r�&�4=���W1Ҡ�o[�&ki�uV��U��S�OO�5?�_p��^7 ~'l��˒�àh�)D�]�98`"9�	N���'��w	�=�X5���8a�|���[iT��!�x˽?~О�"��J�������B瓅`�O[՚>C?��%V�~��ЋT�4q�%�W�ǿC�v�>��8���8I��Sv��������'/�ڪ����e�Wj����F���>���_lGé��z��=dy+�䑹�2���h�jkw)�Ji����.ƒ�#��ch�3���:�:�(��>[��BIN8��h���
fȔ����E����g5����Qu�K5�G�f�r���Q>�� o�7�/�{��`�'ҩ�b+͂&��@v
�Tޮ�[:����Ō�b�R`!��d$Oq����B�pߞ��&��b-JS֖�U�����*V�̊�E�����.�Ղqo�=NLP	���В���x�� )SV�ꜰEx}�+u�ͫ��C4f���?���]b$g�C���(��p`�뒇����rj����s��`۲4��Ih���ٽ�D�F,���p�e �  l&��+���D�F��N8펮L{���J�QXV{8*Wƣ�!�<�@��^���/::��	�,��Ib'|��X��XpW;��aq�1:1��pK��ʂ���U�p�URa6��ۼ��=�5�R[:;r/
�i�!��`�o��Wn���;�qj{+������#�#f�R�|6B
�g���=-s�:7��Ȩ��9B߿��ZcjC_�^\j�q�tR�$>�gA�Sk��}�>8���_�5���*^��zBc8�<K'Q�;R�_���E�vǣ>�A]-g�]Q�LqC��r�.n�xvļ
>�B<�\ě�:Oҕ�6�,@�sTZb:$W�C� s+�����|�U/+��Ϳ��>tȐ��)CuQ�9]���Av0���d y�8)� @H��J$�;m6�kDZ��?\�yK1{z�~�t؄��F�6!�-
��`k��h��M�X����g�H�.B\`v�����Ұ94k>SU��tEEy�l�M�aA�3�)j)�"r�����a�M���h��)�Fʨ��X�[��~����zx ���Zy�Ö�G������+v����̯K1�'��iǲnL�l�I%�P�톧)I�;W.vm�4|�Y�㡊��l��Z����m;�*[���� ���?��A��xh�gxuk�1��U`����]e(;>H��N��׽EJ��}d@���^��Bb���������kK����ëEUH�6k�4h��#�D\��n��[�D-z�:9,.%���)�P�
&ȍ�TXv��',r���QVsn�	q�����xqBs&�^*\�^]����jkZN2y�*�'�CC,�U���a���)mM�e?$<e��P�dqc������]_ Z�q�{�;��މ@��Oڤƿw���Ƭ+���v%���ӑei�9��?�O%���i,OE�X�	ׁ�>I%~�U���"��-DX�H(�hMx]YZ�!��Z A�u{�;Z?��Y����~���J�19��O-5̅��O[c�?.R7j�f¶4�)J�TM��dC�<�i���@���sqi7~L��>�G�v�͡`�f�r�,k�U�D�� ,4�ּt�%�l!b��@�B!X� ټv���pBy�ʍ���%�.� 	�P7'�+&�	�n8&5���>�d����&o"W��K�����_(�9�>)��3p�3��/{���:�k4<x��l,K��F`ͼ���m5���G(ߙ�XӁDO���o�9�4U�0
�@
o_,���,�/���>�������:5�ƍjB���H�sɠ�\�ʗ؝A���l�rQ�ua�O3�wY'n�����ۤ6t������彁n�#4�0��6�04�����1��eP�Ӈ�����T��s�W�4����$@���W��ʙ5Q0��4K����9��1�M�u�)w�.>�$n)jmk�Oͦyc��j9���̃�̮��"8�����u�(�ܳu۫��k��I���ء�M���+�1H�P�2��w��De�t|l��x�2��G�q1� �I��F9H/l`�ɌL���Eѹ�"���~�B̘S�l�DB��D���v��?1���=�/�����x9�LuBG�r<n�8g _�+�d����y�4�i�{�|n9���hs�Ծ�󩫘� ��`��@$��=R�"/N&���!~�8�G](�x.T��|�jI�ހ�*�ѥS��L�{�e��2�~1xeDGº��9}2{������'�˼!�
�H�o�=�n۴��3|�{�D����?[d�?�B�3�����M�S�;iI����h�e�&��+�n-���>y�Ќ�3)�%o�@A�����`���<GhX�G��k��Z�5�؈�����z2�3���Mus!�G)�=!��&#�����J�A��N<q��~��фHST�7D61K���a�b�3kf�"�C�=����X�sm&��Ж8u��0�M�ȏ���p�%`��ȣ�`Ap��~�i���.%�$��7�H��0�=i��'�X$SY�xdG��-櫏?����t��	8��X ��-s�������5�.3mS�n��g��L�vI,l�&*^�ӞE���]�S8uF�{05k��1VY�s�9c�L���m��V�=���9��ڊO�S������ք'8G�ȓ|a�Kڀ�"� $��k���@jv�g�:�d�2��E�Gw�(����
�ؓ����F�A\j�q��a����{�C��BGHc�k�S,����@�p��Z��ua۵W�=n��}�dC�ş�NS���!�lJ��F=unc�Xj�;"#��yȰ������I9ϓ�%b�o%�B.��t�&̅{c�׆Z#�4�:�\���Ǔ�&<��}�1��"#��o����?�?V�W��|��.hZ��~�%��J|$�����
��\^���XMВ���/��Z�y�>��<��b|�7��f��а"����f����o��|�>�M����W�u6� X��t!�h�z}N�8&�_:�R~\m�W=�=l�U�X�X����'-Ew��l|�u�!I������
f\����(�i����c����xQ��Xr��_�Ez�m��0��ǫ10��u{b�~̚2�7����N[H)��]tI�����~z����3��_�����W��Q\e(kP%u���x^8P]�P��q��ӡf^*������@�i��N=����S�ȫ^�F��7���E�B>?���N�4�Έ�@��������m!��:b�\XxJ��/��;ea��Gq�Z�z0����H��#��%X����)���Y�Y�]�>W�h���7���˺���(��<�|���g���ѿqj~��v�l+~=d�!�6���>p�@ۨ�G8��@el��#���S���pߏ�#�3��ג�� ��Ic1�+*)�Z0/�ȡS��oN3�T�{^y���� �+r����F7�����(Q�U�R�W�T���Ѝ?]f�r'��k��sFݣԖh�٪�+�p��T��7���B�(5<)�,�]h�;�k����_<�rO����~i�R:��\z'���0��Lzic�Jp��8-�N丣3wv��b@�%W����%�;�,�A 'G��s��I\�IR���0�p41gQ�AT�7��iP�>�2W1�A��s;���v����6�"�X��`q�T^�μ��?�Ǟ L�vC��|��~��A�@�N�C�d��d]��t �z�晞`����4oȝ��ۋS�ư�L-��Ty>�je�C�p�<���YR�u@=���QR��\���K�~�����Y\E�Z���cGCk�U�=��#��
Ӊد��|=>��s�.�4�(��gc�7��sޓ�rf:;�<�K4<c�L�!��[�X�h>l͓a����p�Dl�P/�(g��rj��~ƙ3���o�*���Z�x��q O\!<��D"DXiH������V�g]/�n�8��v���5pv�H)�y�rЮ1'0(���S�����8��PM�̺EX��������0�횃u�a9:U���TU�z9�R��q% �Ղy�MO	|ڏJl��I7�܌=6���f\|��f76O����1�3Q�
�JX�;*a����A����,�F&���a2��pf��3���P�X������M����ܼ����d��0w)�0fɼ�.&��\�V���f�R~i�E:p�y�.z*�خ��6�|��[�+*G̚�R������3մC݅d�����Tr��u<�Bŉ] Ԗ*͎�i÷0�{�D=(X`4QR�����aD�yv�Y�������y���N��3���g]Q���� O]��FIi��þv��GU��z����}E^Ԡ�M�-�l���e��u D*w��zv�ݒӶ��pZ���k�`n239^���\��ޔe�I'��H���;��	�(��IR�g�����'�;n��hS�]���C�0�iV������У��hT��Ck�֫\�Z�O�6�Ml*��ڡaKC �ZeWȑ-8zv��x��4�1<B;�	hr����0����J9PX��Ţ=�v�-}zhT-���q�܄�߿� �4��@0��X��X��;�\XiuW�R޻�^��\��5���5�����4L,�V��=^�"�==^�����c��,�d��Q�e��(���g?�(~0ӟ�|פ�,sé��7yO�.|_,��l���	�k)' )+�����PԊt��I�g����o��2)������)���jʎ�f���X��56�����4�u��멀���x�:�������0�����~��R.�־M���M�"���w�Ui��Z�̢l`.B��� ��%s-���j0Φ[�m[VU-�H��YF�%#I����1��a"Y!w=���:0���gp��]�o�B����ֽ_cZZ��e�[/���T��E���}��N�	��`���cb�8ixP�)b5� ����^q�fdC�,�O�L>�/���^�>]���;HN�f����ե����R�dA���8�t��s��7y& �K�J����mz�&n�W%�hW�G�h�����	O��Or5��ў�[2,���]�G�O�cqh=7^��e�Ea/�[$��}_�����6�a��g��íȉ����5q����!��z�Ѕ���m8���+°�[ȉ���#�(�}�i��|)�ؕ���R.�ۋ���!�����X���5@�S;����<�ƍ(���H.ɱ�1�Ϥ��㗲|l�����s`��='���"�M�-m�(w����!�����&I3�-�Z�'������P�]g����tgmZ����8*��T����Ҽ��t�~P}&YF��M>u��i�,7���}�s�h�k��Y0��GC��-ΐ����9����d[7P'��3�ܚ���s
D��&eա�'�1|���
O膆=>���B6��Z>l�������>z�A�1�ܥ����pE�����ۉ�oeP���!UU�I��m)\ʴU.egtޗ��K�1��h5�������;���M2}�?��Y`ܛ��π;������,ߩ�7�������mn�n����V	�+Ub�;(w�	*�͋�3�0�!��v��0	�^���D7$�S��X�OMx���<?�T���/Q�م��3����F?kdKAr6�#�!��p�U>r���Z/��;WOҙYV(��� �����XUR�~����QJ���|Bv�+"�o[ ��*u����"iU�q�E�,��a~l�� )ϟ��J��l�}���#�'�Ƈb��/�o��{B 9[�~+�:ۆ�UNPM_?b,UeY�
(����6�2^׎��'��q��9��	���L�d4���F���+��,�Nv��=��Cx���zK~����FocQ���(\/�G���~Y6 �C��G��W1�X#=>bw[�
ŇݚS$���;��D�x���楫�h����u��7 #��K�vw���J��9'U��I:��Ca�b��ݲ��m�6����۝8<TQ8�"�So��i`1Pp��7�^�e�PV�����Q:ba�i�}�d"��(d��&��s�������'�FKY��9��M-ϝ
�ʍ�W��>_^���2y E
�B��!�M�dq���v6!��g��v�C�8dz�X�H�(΋	}4�w����ހ��=��G�Qň.�*A>e���L�f��v���N��ot9uU�v�?:YX��	����d�u��G|�#'�W "�_Is��6�ЩwZI԰H��_�ي&���>I?ǍJn^�\
\�����7����g2;��A�.Vy��b�ѥ�f>a��Ӫ!Ԏ���dΌ�������Ӻ���&;T6���B�;�⭡��1��;��D��zq��n)�7�(�c��hp�K�Ŵ�6Gw�ۮ:��WN�U{)w���r��\�d�.�'�����Z1@���k��.L6��_�7���DOT�m���k�$��y�р�����c���"��LTV�O�Al4�ͼ�`�iMm��/S+�(�����b��у�6�����X#�$p������lI��re1�m,V�ʋ�ںY4I���v��ٻ��������+�Te���D�|�{nk�+ "��H��R�9��k�q�ǡ�~rm(�/���f�>G* �D�����>�x3>�e�3d�����p�]�//U�j��q������� n��uQkG8����7�R&�xs��3����<���edc�vt����u����j����O�9�4�%���	(������C�ع�a�
�e���Ä�?�,�\�O�	��
��1H.x9ڶ2(�7hv�5�pް
J0w�T��P�;<��`���-�$Y�1����-���єȢȋ�襯\$��3ٸ>?Pl��-q�����ҽy�x<�\n; z�݉��V��ّ�z#p�b<�����Y��]0Dw��G�,X�a���{Σ����V1���~�H;�+.����Bx���1�=K�3z>#�h	��ӗ	��WFp�݅@���{�g��ջRcOA��I+9f�?��!�{ Z�,8濕iykg��v+�CN��6i�_7�E�e��:v�����x�P /��(�Q�W�!�.��R\ILoI�Ω�ÔK�Da�>v4��=%��P�}��5�Ȧ+���2{�KZ_�B�}#}rh�	z�t��(|�Ħ�����C-JreCY��0�G@9-y��� x��-� ����9F��Ƭy��oe�!f[�!
����h?�#z�|��)MI�_��[��Fh�m�/�<̇�g	�l��;=�(c:g��M��7�a�n»F/���g�t��1�;�o8w�?3�wC�0�� 0����v�F֪���pʫ�B�S�����>`�]���/2L$	�j\�
����ӈKx�}j�NNN��h��'�a��1g8�5����e�:��]�����B�	4��huF��1J
OU+������^�S����V�R�"���<ӣ,�,�W���y�Pb`�ro���<)v��`	�
���J
�0���r=��&�����;�,ݫIEj��T��\��@x��A�������/(3��Jd`���bi��n�\L�S���	���d8�2[��_W�͖Ǔ=�q*�Qo�`v�����u��^os��#�	�ǝ_��x�t/�
?��T]ZNj}c<{�^��݊�¶Sw��&ڲe�ޕᢙ�0q�I'(�����lrt���6��^�r�a?���ڭ����+Wf��<[$��ܓ�k�t�Qo*ٵ��H��[N��uYk̢�>SL����
PA�2#M�j4�*�>rS?�F�H�P|�������v�5�x�3`>��m$B���*PO
��@f�D�L*�����ݚ}F�#�`(H��kۘ�l�'B ��B�j�ZIk��N"����
^�^Jp�s`��7$��Ur����n�
y��8�Y�ƽ�C��!JdG�`C�`� �����V�l/6�����(	E�?l_	z������,��p�O��S�G>�hM�� �|$� �����<���1_ӯ?� �j^�A�iJO��
`�^�BW�NٺW��}���L�C.�C�c�,�vAl(ϫ�MaV�4�k���a�q�xF@&��+�a�ܡF����Ыe����v^)����+*!o9�n���R4���tk\�ܱ2�s��?+� 	�W@���{���`w�=zf�d�MH�DPP�^f����/�;�0�sV/�!�ȷj��<�t�]��ۨ�L�H���q�Z+,�:xd��
|8��P@��2�Ao�b�@�2�28i'�R�_r�]0���l
$�����/>a��=%�����!"�4�����D����x�(mȺ���۠��tY ��rOj�5'-�~��Ƿ�T=2�mP�>�l�G��c��[r M��q����Cx�k�6K.�d[N��k~�Q�O���LE=��f`kj�>��
�2�g��~M�Y���/���Gzd���8zH��GO3\w+����#
�"�y��'($��K�O���<jb�YH'������.�E@�`����V,I�d���2�o��2��� �̵�さ::�H&�ڸ�Nk`��n���@���|�V��q��jiiO�Cݭ����h\��� �M�G�m�.���X�2�D0�����%���#Q��b?ޣ$|eY���[Fb*�B�h%�DG.����ph���g�����Xkh?� �Ts����t8@�J�;��6���%�o��3҈����u�:  9��Bw��Q�P�;�g1t>Ji�-ߡ��8�92�G�桑�5�+d���	<mϚ�����s@8���r}��pǋ���(a9@w>Om��q�Ҍ����[�ۇ�.�����<��S�o���=s�����C�ύ��$�Ucw��s&t�kw��,�h5H����Z�^�s�G*�@���az<(��?�v*�)�1*��y9bhp��d��'�H�9X=�-/]�D\��d�~�3�]О�B�SR9�n�-%���[Q�.�W7#	z�`�M�������������]E��[��)=U�F���5�^��c��Y��� �Jݧ������g��/����Ӣ�^���� �����n�X�QLߨ~UD="�ݔ5��_��B��Ư��Te	yI=5�c����Nx��a��P��q�'7�3�W.���53�]Y�ӥ��s���*�Ϭ�jK&hvb;7��0
k���I	��E�7s���+��X�kld�{��q�(�	����g8�k�|�)��;�KX(��ɑ<6C����0�!՘��gg#tƭz�\b kO!1W�FƤg�z�'����?0������hJ�D��k1;k鶲�(c.rx�_�5^�=�k��xz��50����O=*���n����M|��ux]|E���+X����w(Ԧ!5, #+���H)=#�����5�xR�k"����ɯXȷ����=Wy��k����ʋo�:g~�T�W>�����������Rs_Ҵ]������fS,	n�1��jȌ��`�sp�/YƋ0��H��L�q��\�*�
3��:[��A���vJu��ӯ[JMx��X.h�ςٖ;�>�-J-��W~�"TOd�cI�R՟9���kś�-��v��p�#��	��>b;pF�i�A�.I�*�4�g��Si����l�b�f�,�]��H5�L�w�L�]�c��@t��<�������%�R���"�2_�ߛ�:�$�9ץ�UIuA|��ք$-b���m�V*̈=�2�/�V�g��_�8=���
#��pJh�;��3�>����9)�Fp�Ƞ�+V3�+����p�=��	���"�`�����Ùu5(����Q�kxI��q�n�D�Aյ�CDۛ��L:)@Õ�,�ӍxV����G߫Ǘ�z�@��-��� �lU'6&~@�6#ҭ8
y���u]Lry���S�s��������ZE�UN����
yn��(Z��`���W��a�'f�j�C+0�[��P1���$��A�{�h�bcU��K�������5r�+	�9�|,i��LOeK��}��M���Oe*�mq&��>	m#�:�"��Ѣ����
�Y��N���2"��w`�'82�"��m�W܂��"�}>�- vC3�9f
4��cxZt��,��E�V0�Ǳ-	߾�9�/l��ϩg$a�yڃ��(���b��P���t���)����`h�_$�kVF7.��Y_��81���c%#΅����,7����?d�������\U�M&[��7'j���6߮/q��+�(@-H�[O��C�^t�c���Ӄ�7��u��AM���,$4��༩��Ѣ�x��>���^)R,��0�F�ΤH�lT&@�k\�G�L�$%SV��b��e��Kxŋ>�=�tJ]z���I�;��-޵o_Y�%U�5�❾D��)�oȥ�|����`��d!!2�`,%�96�u�4A�oq0�9���b��nF��M'�HF�KE e�H6�!3�tV�z��#�.�����L�'])�N�)=�[�d}��`�
*�.iܺ���fG�
�� '7����r�l#��x���oO7�|]4_y���5c?���W�=�e'G�Rv�A}��
R�+�g��I�n��#���8��Q�.Cg�6D�3�
s.�;+d�:�B@V��d�$�%�3��:N
�^D-���4�pؐ��rh_��N�}x�l�Cf��h����,� ��ЭD[,�Jr�ⴰ(o��M�}��8�De����I�W�Ӑ}�724� ��o^,��֙C���_@�>s�y���m�����s@�PY��Q��P����I�R�5~�^�)!W��tV���$��x��1u�2�}�����T3�����x�w|�4�6�VΥ�AF�
s�,��V
���>�Q�>�gd��^6e��%w<ZS�M���9ߪ⊋�t�+� bhŬ�ZɚY���X;�Q���^���D�6��_*�sd��²o���A�P��}`��(�;��y�jmY�����SFc�:L�C̲\��ȇ{酆�i 3�M��+�Q�ӦP�
�~|��W�My�� ��%,��
�]��OI�s�ZQn�i���3��F��2J��@쒈���:�
��ZǠ%,�����YDG�ڜ��/r;�GR�>O߈SY;�\T-$5��s�����Q��Zm a��g:w�%���p��OMqk�O�&SB���7��;��
�b�>�:g#!Tɢ!�d�=�]�]�������O�KO3���P�������i��e�F���Fky��������-awp$�PS���Dٖ���{���@|_հjs�,/j�i���`�s=ִ�e�����D�	vW����=��Z)y�痖�	�<�O�T����i�JCI���N��^�yt/y'F����l1�Nm�㐱�GpXȎՑ�&'cl��Owp��F�Y�o&#Ԉ_ˋ�Z�Z���j,��b C�U�к���+��Z�^�uHK�lm �rcF7���uAk�-<�ef���Kg��u������3섷��Qn�e+�:�.�:�0��n?h(l�G.�-�i^ðBD6�$P�V�!m����~J��ː��7Ɛy��锘
�)�(�I� Qp��H6��k���S�u���)������3��m���lX�Bt�mH�\��FSi�,���F#��kex#���;�r��>�G.n�}Eo}��}�� ���)���>��~�xq^3 Mp�Z����vf�$�w�P̹�.xe�tS;��m5/*k�*�J��[\t�m��>p%�9�j{�����	�p��3_�ƕ�fǮ��${l齬t�r�G����	�G8�#w�h�k��43���q�����ٔ���N�6J(��\�:�����(�)
�Յ�Z�zv�|�U��\q��"��,}�����l:�26��8�,�NP�vP�����]P�/�o��#ᆔ?H=ن��b� ����%$���(��i �:��Λ�+{B\&%b�tk��&�{Nr9�w����tB�_h�.4.�f�,{V�r�n�jŪ[���-ω(X��9�'��latñ�!�U2����E�-�����d�ק�჊t�0_�A9�U���$ٖ�-:&`���'�ob& ��Ku��(��	<)����8"JV�ۂ�k�=�ѿZ��J2O74��l��2X>g�к�w6D�e�+��U-������:���B�& �I�\];�o�4mPߗ[b�����he�0v��.M�,]�J�^�q0��qSCo�M���*�6@�2H�Vp���3>�#��ٻ������T�{�.�����lz�ې�h%���s�5�|0
���4P)�1a��J�"rt�"O���]�y�6Ȩ٩�`_F�2w���bN�OR8��S-.,
%!	)` .1�s�~�]Y\/W����3���fI3a�ZQ�.$��,6x �f�Z��=Q�OJ04����^o��[����eV(?��,��Q�u	d�"UI+I� ��e�$O����9q���d�4�� �����S���kX�u����'��[5�X�7��r��!��8���+K��f�OՄ���
�a�%���8��W& �����)��8�4n���ǅ�5#t��E���E�~s��5DR�	�23x����ܣ��Xm�L<z�����#\pzT蓜���%#�`5.�c굎Ӵ� X�[��٣d}��g�%��x��69:���v�>	=���
�\�Y�?Ɲ�0���(]#�ޝ���ۯJg:��^Õ9Ghc�x}x��W�z_N���~����}�����dMyW>���¶�M��Q��4�Ml�n:(�bx�s���1�r���i�Z�]/�iO�W3o���F�<���j!����;<s?}'|�InpT)�����/x��K�Ŕ࿪[3�p(�j]�HP@�g26��j��"���^WH	��~����z��؄|t�b���B�K�}߽p8�be�>�r\�b�i�C�Q>�J�U~��Z�kV�ۺ�nB:k5�o�K-����8+V���	29�RL<W�d&�DS���6���Bܜ#d��DymkqZ��
#��;Gg</�˜ͦ&��)����8quM�x9fN�ږ�5ʅ�͎E����;q�w��g�6�3x�|����[��j��>�<0)8��;f�0c����kzzӛ��+Q=��y/Y�N3�[�G��"���-��^�n�r��)«�}r�<�K�2�	(ԧڑ��"[Ċa�믦���c�T�6��w�Reb/Qs(��A��jMg�]s���*�$5r�'u�*@������,�em���U� �ދa����3}��K�x3�4i>qo�iMP�9�c	��-�jj=����W3Ԕ������^� ���i�jυ:]�&u�Y3!��֯t��$�&b������>�;FȬ�8�?�}�ѵ�X�T�Df>D
<��7"�D�nC�� �q�o
rW��}["Gu�厾²�C}��H�,e>%��$M�qL�O�$_��MM�?�U��w$�[xDf>��SLIn��+��j��o�O�����*���:_)��L��$dW�3%�8��4�Q^��6�Cɼ�w������j���'{8�Ԯ]`�x��F%��2a0�b���xY�ć)�����$F����zx[E�棾�jթ���5�K�BH��!=uU�$B��=M�� ���Y��]���6���N�=}�l�_%Sc���x��X:����q H�aH�|Y�2ʉ���п�[�R�~����l�����
�~(�$٨9R�z��-�H8�b���᭧�����3�E�C�T%d�?�9�@p?�Ȅ�p�``�+�pc\��g��}�	f��߾��Q]_��E������j�N��v���Չ�XV��*(�7�=a�^���>���S���4R�3�����}
��^"�CS��Hұ4�%�kW�.�8��ь�K?b���e