��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V����hN=��a���)�硹<H��׮��`̼��D�g�;�mR�#rj��S��k@'�q�/�ha��pc�R�(��g�F�ו�����`d%D��G�qK�DW�+X���iv�O�O����9�t�0���`�<�F�2MGJ�g_Ю3����Na/��4-^}��ru1������>�9��& c�dN���(�lE#���{��5�h�ɉ^�F8���>�%8�
��=�v�����6%ȗ#lM��98H~�h�Q]f�����-nf2}$(����3k��b&JX��8c��ܜF}H��ti�;�?����se<~k��]���A�NQo�1����~�t���ϒv���B��y��5JZ7�w�r^|�a���KW�yW��5�G�ԣ5��N����E ʼ�����N|ߩ��5������l��Ѵ����|��s-O	�>��7|�MJF�q�x�:��)��KQ��a���
K���}+�p����+1��JUܢ��P�<y\�
�~9]���I.�6;t�O�nӋr���>ߜ�X�2+ J}�5���?��ݠ������p+�w�>Ѵ
�>m Vپ u����f�9��a;���u��a;z�� O�����[u�� &jư�	�=>�H���kfj�V+�e��Ӈ�������[�T\��� ��Yx�)� �z
:z��H���ٶ}���'�'J��!�:xb��H�v${���}s��������`�� O�t�|I���G��C���^�M�A04:K���ŝ�Hcj�9��[����'5]!10�\!�;pt�T�~�#iYy�)����V����[+�=ƘoZ���>���I~�T� K������-R�}o�8�!��m��AD�ىPy��R-X7��#�&�|��"�����ǧJ×}�;��JnND�]^Ѥ��i7/B���M�r$҅ ��'2���O�х�[�A��/�5/y��P-v��'R`It�v����K#Z�o{������bI��5� �^�Gr�F"���]�͉�@⡴H��w��=}�#�~|t$B��)$����݇�q�C=��gɗ�^�r�Zo���ܱ7��
6��!9-�O�%��C�C��	}p��f�^)�E���L8�^��Qy�Xޢ�,�
�W����A�n��Eg��#t��_�J�
r�X������i��ܟ,3o��KOJ�FL��	dVM�=%��Ʒϟ�j�6>N���t��	��Ymx�_��M/�}Mh�^H��f�6^���!o=c�;�$���p9bZr]:/��7pJQA�X�������)V_�WE�:7A]��L�����/�ƆoA�ۭ*��w|<���*4�0'�;#3A���}���GG�n����sìC���iL�y8�a��L�A�G���:�FC\S�f$�H���h�V�N@t���(M�9��w��(��o���ҝ˪V�|�(}���fH4�)
�����@k.��7�CN�ϖ`8#��]C���<��c�ݦ�ۊ<O�I���Y���� <����xж���
0m���P(�.�c0��^����]�]���ɷ��͊�l�%ՈUQjp&�Z3�'�T	����}�K�]4�FR%����J�X]L)IE�)w�םQ�i��a�?)�����d�#�1�2�?c Jq[�/_�y��.l�Z�� cI�+��jf�S� n�Jw���<9�r��~�'r�1��,����U����u!C�Y?�v*5�}�+G�R��TJ9|ϴ}U��ce��Ѡ���#<i�tΜ��%�)(0��l,�BlK��t���CZ�>S1��s`��'�ur@���@�kJ�"_f�0�%��%u�c�4�[H3�Z�H�:�j��a�އ�4�:>[��/�^�S��߇�(����brO5
e�0?���E��%�z��� ��IrhI;�s# ��>�e��0$��{��΄�m�R�����T+�/�&����a�r}�q�\����aJ���0ogR�^?Q7f���&�0�l�[�� '�N�䔍� \-!���9d���|�ʯ}�IwJ������?@���4�f�m�n�I�霫{�0�4�<h��):c��:4UV����m���tGf������C��µ��cTn>Hk���z�U�@ �Z~��^4��&�1�%��ҕ7���`]�|���	�wVjnw��;�f~1N~
O�.�E����� ��b5�]��J�o�~E?d��)t�~11c��w�*��O_���: ~8�{T~V?�Л�!�?i�ŽW>�7��!B�S�1�xM�i��\l�`BVjҪ֫����V�5y�φM�,���%�*�71����WɅ�Yb�#��`��X��C�����ڀHA4�����V�
�%k-�hz{�y&�^A�d�lS"�]�/+���K������c]��#�2'[i�W4DU��׳Ŏy��	����2��@��i@">��_��-|�-i���=(�CJ+���C�UTGW˨Q��4b۹j�"�|���7����B��0�	��kF����Ъ�v�p�-�X�|�h*�ibܔ��2(�x|�V�5���p�{YN�N��[}���5��Zz`��6�|as��rp�� ;O�
b��"S��}*6�wH����j�'C��Xɫ���H#�Z�ߓ��ri�ù���.o��i����#��rѤ^"�]Q*�s���W-��\��~Xp[t��3.�����"0����V�#�Qu)�	�C��*����[t�Ec�6��\�NN}��m����C��!���-Q�t�P�����-���U�Ӈ�&Fpؽ>�yոt]˸c`	/d�@��]���Q&��ձ]�@%0�OKg��mnKz��tI��PE2�G@L�Z�����-���8p��)��b��6d����i\���JA�x��K	�O�=�F�?�R�\�8`�we�I8Βn���z�Tj��N����٩��S@o-�	��q�j g�Š\���l�M����kY��+�Hrک4ʠ����$�X�R
C�- z����L��ziL,��d�Qq��_��n�Pŉ��R��.���ppf9��A�Dۑ�K����6X$��m�g��D :}�>.��4���R��X�<��{nd-���9Q8��f��g�>RcV�������4	���x��EU��2�M`Ž����ق�r�"]�2�P#��(�׋��ݫ�Ci�vҾ�,�_~Y bZ���ۘ��ʊ�	K'A���RY�Ps���O����vF̪>/�k�`�KeM1k�JIK�q�� ���b��ʚ���O�F%tZ���{q>�XB�Ï�l��f8��cW������lx�ێt!#����0���ʑ���4~����S���'��"���y�u�������_l�q�^%"@R�d�k��ai<�Y6~�NC)�.��9WA�C����[ʎ�=sӆ}1	�E�/Bt�ׄZ��Ԛ}�0 �YK�������%��P���b�Lu2w��0;u?G3/��ns��"h��hL㝔�ct���0�:22.�X���/���<g�+�\V_fUamВ�,�+]���Ӄz��~�K2m����:g�n jx��e>~��|�\��B�Jz0���䴰��Kk%ֱޛ��(�P��^=�n=NZ/�*���o��8m��	�<+c�W�����)�#�&�t�d��K�?
�d�&� }����,K B���ȠZM�Z��-p��O�~-�9jPT+<�e�Sl�}O�K���m�e���`��g��Wč(70��u��
�m����� e$/��j ����κdnX��̓ࣵ�3\�j���G��O=�Ǎn.���}��mv�[�Ҹ<�����X����J���[O�:�Tmt*rBYHD�+/��T&^ wn�UM �I�T�s���+�<#�BR�ʧ��"�,�mS�]��T��~��Ao��9��K��f
��ˊ7P�y~*��g�>}�Kݓc=�8yeg����H��x�f�R�X�^�����>��K3R����r���Oq���ՙ�ׄn�%A��Ҭ�3�,��!���Ch�s�m��7�\�2w��K!��0���?��+�������3����$��_�XLh��a���TSI���r�>��1�����-�&2�ʂD.L/b����fG�M��7U���|���u�Cz�	��2T�'o�ȔU9�9�$�c5h��r�浔T�7�C����>���!dYW�����{�Vwⅷ<�0���hd\�vl9�Y�e�i�1�b7�uB�V������q4X'?b��7�*,4h���X�j�IY�l�5����4��vAl �jm�A�X�˲ؠ� �y��d�����b�R��I���(wӸ�)�]ҙ�ʜ�{n��T�HV�cǻm�4���	������[bH�K�⩃�嫉8���>4�$����0�Ć� �ǅ��3%�懍�U��&�|�q\�0�j(f`��U�Itn~�.iz�
�5VI�����|��S�s�/�6��c����u�w�'��R�_�S!Β'���R�) �1O|��N�WED���=�P�����L�ԡ�z{�f������~9Y�i���\�_q;.�'ԪDطhv 9aņ�1� 8�ޅ}�`A�~�i���E�����q@�#8.� ���{��ga^^�&˧__���deC�=�nT��2�/U�c��a�|��9�G���S�9�Lߌ�;��&a���^U���*Z,ag���ӂ�}vot��p3��<���4��k���3�ޥ&/ďH���
nضQ�AGP�Qz%bM��R@�-{�ܻi��b��sJ��q�>�ШA�&�U�<��ɿ���j���Ѡ3jy��m&t����*��,{_b�k��[5I���UA���L� �w8l�I��m��OfF�Ȇ5��p�:ht���]Է���7XU�-��O��4�Qq>��G�_wh���d�>�p��0��tա����T�I2�ƭE1��#�2�G�/������Wz�6[2�c<C~U�	fR��Z�z��8��t�����-�v���Kh ����"��X"���r2={�I��{�~3��K��B�ϊ�� �]��-�ˮ�c�s~*t</������%j��9)�'��ٷ��w~��v}ħ�V�ȏUT@�L"%�����M�n|�2�� ��kA����>�g��� Y$��Y�U�"�p��Zi��.f3Q�#����7������ܣtt����ʹ�7+����de������̲����7����zݏ74;�ۀ�!�B�.�q�N�/�9�NdSo���`�\�˫�mC��a\.�n�^�V��wC���u�!�0W��K�L=K#,��s���_�v��� ���#)�t[>��46*�C����r��S��V����iRZ�*s`�}뿣�2���Ħ^�����t������ݜ�G�;7yE˫7ٍSf�h�U-|�)_+^��C�Vk*2��!NSz^Fe�=����ώ��Nd83��"�xn`�:E�H��M�yx|\k����L\vK̦gx]C������?�$�P;���e;N�0�iՄ�4�̖D��Ʉ��H�/�� ]��dk���h����r��~�ܤ+T��]�}Wt�e��*���M�)�I0���>"�7ښ�P���v����7x�c9�C�TbR��ҶG���1�:�=7mq\�q59�-X�p�f�ےx�^g���V����O�-B�m^�$��wx*��uV�M�116��Cr��*�^���ahHE%�����Ĳ,���Q!�Ea��,N��Q�+��/%�y�G�X��=��
����Y���Ch���l��p��T"��izꋰ�U}��:+5K�ࢯ�aQ��f	g��̨��SO���f7��AN؀P�2n��3�ב��b�r�z��(	�!Z�����e �������So`1�Sy�${�G�0nZz� t�\��ݘ�v��T`{��,u�v� �V�]���5�k6����-�>�=B�	 �[/�R^q
�>k�o4�kr�ϸVM�=��W-mM�,Krq. Pw$�WWj�`�7��TU���͌�Y%C[��Y����0��%��,֏��vI��8k��/t������_�.|j�),��rV��n&���`���Qf�߬��u���1>���:��&O{r(��2�h���8d(_����aF�م�1m�f��vQ5 $�SD[O�Ҽ:o%�$�e�mIYY+�k� �{o�~��-_������I��|\?����A��T����YI��o���|��AL᳴�w+�v�۾���K7T >s��|?Z�4�O!<>�#E��kH����.58�#��Ad��Q����v�CX�(Q�J2���37�L3�]P�R�'s��s�!|��D9($�f“��2
O��(�c,���%p\f}0��MT���7�y�o�pM��&�����!�@�K�zj�f��9��G�� ;�᭛�%e��x��s0h#�[��"�>��;�i��#\ ���^����l���;A�D2L�,�jd�oa�+8��↑�Ď�)a��ba?.��[�bNkt\�0�`�Jض�2����3�|s�@�YL�I�}c�PF}<;\��S�+�	]뽼�U$O��E��G8�hV'�x������CV�]��#6r�OpjΣ�Q%������4c(�Q���C�Z�"ļ�r�ݍF�m`�e�g:`�T��kX�f��bL��[�,|��0�[MG!T\:t��a��L33z�:�;C�q����'�n���W��	�: �������©K�f�2}��}��)I�1�۴';{����H��ł���Xc��C�@y�!M��Qv���&����*�S5A��*�Gp����󏡭��˨���[6��{Ld�L��#���4�h��|�CD��l��-	*�G�V�cp�Q7��A૵��:Hm�akl�W̉"�����?�|Of}��� �o���0(x��; :>�%���۱�'�����/��oy)��p�7ڧ��½��)/O�1(@��w�ƙeҢ�\t�f���e��FKr:ބ?d���H�g�c[ӽ�=kK�|tz��m�lO7��:�3�h:E�����rH�͟|3G��N-��,#���u�3��gA�x�c@�@���E�/Y�L�r�Jg�U'�ݪ�$O^��g�l\��k��Ճ6�E���/2RFN��$���PG6p��l�� �팶A/T��0n���Wa C$x�n�6x�~�f�~4�_����W�"�eտ�q|�mG�3�H	�U��>��SQI�>�!Ϊp��[ucS4Ee�Aw�6k��$� h�����Iԧ(X�;��r�n�_�6�l��~��(hw�Z<-�Bä����o5rZ��aco�xS-���.�.y�8������{Fa�D�u���1��#Ӎ׼O�^��Dl21N2C��A��(�.C��m��oW�x3]��3�Fႉآ�t�d��|���;��j�$`O��
E@�W {hȾhR�t�֡em:u����Z|9�#��4�[8��t�t�bE��	5:�!�����pQ:s�'�|���:#�>x�S���%�7��>AF��]%s>076FR�Wn�셍�Lv+���>ĝ_~[��km�j^]���*�a�1�t'֓�~D��[���љ 19����4�1��:�|Q#$��m��}1(Ò2��P� .W��������S���Zt�tTHR�"�b/��|tf�p��Y!��C�KK���
�X���4�u�Ӹ4eN�����М����.�ꫩ�,u��X���a3Q�T:����sYm/�t�*�K��
С���=��!慤�vI�?L) ������d5��1�z�ț�Ӗ-�Y�(`��p�(r��1���� ��ep���"W10EoKP�B�����y��;�_��!\sjNE����$04G^��0BDV�{.��7꣨!��O�IY�}�9�m�������\�����9�-&E��!*(}HňU v�y�7�xȜ;�(��1��g��-��*i��1�S�E��I`�~D���$���2���̨��<6�R<Ɋ���z�jjH$�#5�a�J�H:p��l���Tw��Y2����ʓ�ϭƇx��F��� o�Ln&���>X�.1}�U����N׮~
enQ�8���t'D:a3�]L���]+��>�L��{��Cn���Ɓ�n*&�rlQ�}�x����8�1����eQ�Kz�꾦��K�d�P����-��謁;,�6<�ܛ���I��u��9�唁ky*�k��Ɠ.)h�[r
X���]Ԕ�z���,YW~�Vt ��<�4���|q-̽w��7�c�&o����Y�AZG*�'��7��C[p�ˈO:�*/
�)L��P��z�h�znǨ"�O�t����z�����5���(��{:�t;b�U_	���'H	8�OU�{��I&}7���G�j�3�?2��J�5�,�ԉ!r+U��g��sm������	��)}�[ �ۖ�:y|��ͯ�R�W�{{�G�3R5L�!�D1b��Vt�$���48�����[��cJ����ZQ
�_:iT5z�+��Ư�E�����<��\"eb��������%;2�����ݹ�b$�"�7�V4Cs��M
i�)L�����Ĥ��!vɡ+�B� +���W�'���Rx(�G�V2��AŃ�B�,^��l�j���i2� �{�l��a�L���K1�8�f�I��e�z�m���1�ћlU�&)����UmP�`�K�ž�1;W+5��v�<9!�ꊺ��.�q����b	x	��#�d����A|���Z�z�[�C2�T^|�ttB{��<��?�E���P��#���޲��Q�r$:��|{�Ńr��uf��	3 �c W������+!Y(����:.[�h��ޚ�����7�0�7x���l�m5+":��1�h:x�; Rxn�n�e�ĥH�2DU [��X�E��E��a���/6�A��Z��,<���L�Ax[@�F��:`�`r����l��1Ԝy��^N0�̕A<n��CY��mk�|Y����h6r����>�@�B�<Hf��_����y�62�_���?���C�G31;��E��RߚR���W+Yʗ,앿r�9)�C&�y-N���|�2y6l�"w�zg{ߕ���αT�޽�,|�ɗr���_ԉp<��>ao�h/�Y����G��Հ�{�`D���?���mĦU�(�W_�d�('_f�cW�1v�xJ/Jb�#�������}N0M&/Y�������d���;�{f������{*pGۂ�Z=��A*�?��{��+ȑ�+4ƀ�IY����ꄫ���g7�ܩ� +ư�P�i�h�!��R?��p�o�ՋY��C�>YY�\�$6����.H�*b��T�G9 E��(�~<�y36���ٽ5������H�I5�:aʧ����z-��.��,�T��	���L�.\���9CC�K�jy����2{���B���3 
��!��Jl�q�]�g����r�b'�~Ҽ���i��
�{M��mo��q+��l��co�;�j��C��qT���P E��>.��&��T b%
 �W֔�8;"9��P��V/ �T��9�n*����6����d�:3��O-�Pm]��@'�=Κ�<�ig	meHr�)�7�
�F���+g�b�8wR�b��nv�� ���#*uZ�B�i7Iф���Q��J�V�d�$��j#Xo���mB��hSZc��}~h���,܄s����d��T9y�.�y*�fv ��o+�.
#Ly.
�mF;z�����w���"ȹ�d�C��Wj�s�94��鵑˵��F�1vJӽ`D(�]D�m
�^j��6�_6~H(�9��F[�"f�:ow�� <�h��9�$����x
o����6��eI����463Vb�V�3�����֐�Nxk���������� Ī��	���a�I��a{	�X(�Rxec
o�n�PT�"5�ӳ�uqr���FI�>�s�-���_�PE�+%��:����T����x��s����=.Y���F!�=g9:��@�O��O�Me&V\aT��W̢���3�鲾��T2�p�"�ʷ����M����m^�a�����R��fZ.n�$?J�~8��ϣ1�BP�����ֵ?�Hd�&k�5�_����M��䧰|�:���a5p���Y�9�L��������"��L�u���@�)5��#��c������
p��N̷es,bv�>�ť3'�����gNR���٢Ҝ|=r�$��	�2���=�6Z}bx;���p}bR���
 YU�n$���#�W/%�;آ�禷�*�B�BC^YP�R��C���.�ŷZW��-��#�T]R�O��(
F	]3��\&��Ļ�=>�O��{���|���0�X��v��:�t�w#
�"�4z�����{��{Y��k�{��mc�/���3y�;�D�ۭ1��L�~tcK��-�Ci��w1��W����ݱO�V�Dض���s�4�M���`�fN� hw�I��ѭ��Ǉl�����j���` �*A�7����z� F��	F��f�N�L
u�.���9`P*���1�Z,���ۚ�/.ybhFic�Z��@�2��?&�]Q�4��G��@�˼ȕ��@J�`�+�ć;%�%���|}�N�MW��5my��p��Қ��r�Pv{�A�c�g�'*e����#"����/�n��ot�KVA�)�&�2��?�o�_]����f�N-�v=���/��|Mqz=|�0����R��¼m��T�̀�LMyom<z�JV�g�R�5a!f�,/��5v]��Ւ��-�]��f��l�`�7���z�	^�z���EO!Ȫى�>��� [B�էG`�k�"4%�y���N��bG"Q�S�쒿~����h	> �!n�l��1�q�\ѡ�PL婰����W�&R�f9Hn��|g�Z��ఔRM�W������R��a��>v��f�#��-S�A�ל����t�k�{�ђ4~� $�