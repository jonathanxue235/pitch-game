��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@��D�����{�����}��Ț�����@u��=ȳ�V1�RR��gt#qYUX��̮]��"T���bQ�i��������!A7</?� ٘+��)��`��[�^g=z4������Nd��5��/Ħ-�]^�|2L�ݵߒ��P62r��e9��]���E�2��yH����}�2D�Pn�T,����KW�X�.�a�A����a�+�;����$�Q��ȋ�AA]�7��5R�⠳�� �M�Z> zU�d;vZ��>��	��A�ȿՍ'�^�8#��w�����[Ö^o,�}��<�cƴ"�2d��>��3�Ƶ�)YV��2���	�$9y�J��z��/>*��pi��هT�
�<Jm]�ׄ<=��s�B��k��Hfd��B���κ�9�	sA�W�d7��0�����9�(���Xx��L�y�e%%���S�L�N){M�dY%Kz���C6�/��7o�����@�n��h�˕ꭀ�C��@��Y��� ���?�n;ޜ��a�� ���}O������`�Gi�kߌ�X;F�`uG���֖��Df+n%!��3=�ē�/��ALv��%V�����t���RN��Eu!a!�^iyRbe�r5�-v�k�W@�"a�5��>ÕLS
������5�Ȣ.�V�3&�Z��)C�>��/��F��*ѪB�q���#��H�ID�7���$ٻ�UB5r��~�Ʃ�Y��$}�b���Lp���A[P-�{tΎW}2��o�RA���&����h��a��|r�j��rx�AQ�&�H��F�q�(ޏ�a�K�fv�d������������4-1��vɣ�e:PSo��+�fW-�O �0J�&AY�`�N�����B��w��o{\y[!-�ZC9���~��{��|�G���5�[iN�Mg_��sL
�H�����Cٞ\b+�`P����>��Sߧ��6�?<;)b��d��ht,JT�����5���#�C���+>�����Q�?l��#��%�a'��YTo��q�%#&;��; ��ZN^E��`y��Q�R��F3��Ma<�6&g�ɹ�Ɍ��A>��?�`��.{�8.��=iY�d�\?���e+I	����OE�P�`�^ ���5�j�+uvw�oJ�WI`��_���{Y����6���r�+Y������r���IP�
N����a��䂩G�p'��d����K"�s�����\Q�(��xo�H�[ �Bݓ	�g�n#�]{Щ%�rq�Ӫ�[�>.L��^�ۜ�&��� ��;�羽p�湈�G��ᑗ�*��3/�U��e�M,�ܸ�=�+[��^}N��5U_���sގ�ӬΟ��T͢T'��i<-��ȋ�eܭ�Q8�_&�,���}9���;�/��#�C�qA��n�(l��H[d����.�����d�3�D'M/*�<�i9w��=�i\v�U{M��h��H�lR�? ���Z�p��3(��o[L��� �ڵ��O�7��6�
un�t��������1jx�-	�pC�����A�������	Gn��:u��&ԋ���(�WR�k�n�cռ��܏;6[0�g�v��X'���i$�D.Ԃ�4S�K@�G�w[t���?n���ii����|l��ԥ�M�$%�gCc ���m@�k��YX!��R�]�ib��i������P���`��=-�<������"vL(��s�����>��4C��|h�ᖩ#�ֱ]���򿖡z��_�+�K��L�S��6�D'C�r}�?v�� v�TI����4P�3�۠��8v-��/n��l�|x�Vٍ[@&7y��_ZdT��a	��/X#?%3�n0�4P���EV�s��D�	+�~�L��$��������f�\^]�y^��U8W��I��'ᦰ��\|�:*jG�7/�Jۍ�'�n.��8qD�#�%��S#�Hk8p���\5H,1ͼ����`?p�F�TM�����Z��ס�z�����_3�g���w�R�r�
MAj�`3�j6;��9-��,b�dB�C/w]��V����1L�*pP}�H���$����

8�>�!ϤO�ӰаS-"C4�l?���{M58_�@i��X�#��ga�C�FH}�	vΡ}�Jh�=MK�g�wF�c�]O�Ae˨�`@�r�s�u��l��Ɨ���"��)4K�W�DM���ֿ���w6!۾�n�ebZAy���ug�w��b�# ��z���<|�����Z~�b��I��ƞ3V��@yY��/����(����l�V�熖���
:�UF�nP|���akH��v�1�",��z\�.7
�	>=���tw�{��2Q�Ț��������� mN�;([L-:yI�_�8)&j��?[�4���Œa�y˟��`�d(�wן���5}��a�|��Y��jX�{S:��������"w�ޥ�D�>o��y�*ݯ���ؾ��"�G�j˿0F�3?�����52[+#uO�jD�����S2���i�$�%�7Z�ޮ��;����?��"i����`�8�5�n���s�^��r�|�ن�T���"�ɼ�.�XG[Y*�!og�%�!���k\B��	���6�:�L�@�qJ�)?�c|-&�.`��`��/��HH��UA_�L�����M�3�=>{�����C��-�'���
���h�d39V;zp�m��h@�:�j|I�)a�'[�<�b�k$;@�ϣG�G�2`���kC�ͅ�8���eD�c�`�U�|,���O+��E|G	5��f��z�q��f�]P���k�~1��zyZ0�/9O�e� 5Hۧ�#��g�
�0-��I����V��)�O����{���i�\v|�N�֖*Q�$��lt�Ef2����n�"hu�-��gn��w�5q*��$+���۱�x3�ՏPun{_�**��ٴ�v�K�M������}������(��q#x���M�Wwu�� ��'�`�~B���N�tJ��r��jg�F�Œ�X�6$Ž��7WOɜ��sI���-����v���e���qUy���g�ޓq�t�N6��b�06�_��b�~Wo�͔M���z%����>�;�QH<E
!?�w��g �[�����`IT[�^X���<�E'������w��L�{y�lC(�8�����P�߈�#>s�DGY
�<���;E�<�7��d�E��f>�ڱǹ��e����-s*��~˷S�pj�y���M��C)����1[�xP�h���$%��E��k8��8�~�m�o���>���Q��)`�)���ZN���Z��_'�q_/�̄�X�p��66�M��D];�~���: �!=�\�H�ґ�u>Á/#H��aՒ�C�:�"T�t~f8ʏ\�3��.�,���%�4�}=��#����V��%���T��.�!�=+���9;Ga��yx��Yt?����oO
qz�S�5Y�\V�&�̹K��O�c��.n�*6�<�`u)��;��fcjV�������Mg�L򩤃�����J�TwE�L��׹�M���y6ұ�O����`���a�E�����i�!�J����"�6E��F��Pv�ej��|5%0K�~��bk�k7wi���粽mz��hoJe�gK� l�������C���>�Wg����Pjv�x�0 ������@���f���*��L�z]���
,�n�>x.��Z�Q�P[�T�~c�EV5�ܭp�w� �79#�/x���&��e�S���������N eT���ߺ��#��<]���Q�ޭpq!H\0ײ�i��ي6�����O�H���2-�` ���̊|��Y��B�ɒ�u��np�z�
�{1J~��f��Y2"�>�U�<'���i�1��.-
���	J���ٻ`ّ���j&���_sh��b���s[F/����x:���:f^�D�4��X��Y�Z�9E+n!j���t�PfO;p�@T�]����G�+�����{�3�C��	��Z:ɾ�z䖨�JR9�	��X��^��y����q��D��tQPI�6S��U��[|�x���Y|�����m���*e��)���^ޯ����?p�?��秿,�3����OÿV�.�% .	'm��a�+%q�|��}�0"2�so����T����i�z��9M�oO�åvY���&��3�d�Kd����r�'��d$��Eu�];�R�O6u�u��Rm�@)���XHT1m�?
�7�!�#�JY��q$�L9ڬ:�ӳ�Yz��Ùԧ:0t��l��������������HW��>�)��-��t�ʦ��~v@LI�|�5A>+�ayy�U��g���5<W_����J��ǈ��풰�L�.q҈&0��>������I�������Y����!�
�">(g�Ǝv��,��ҷ�}����?!*�di�}�l!f/��h��V�� nX�[WbǱ�vA�S�ΟN'kCi�q��x����8�>vV|b+c4SC�4Q��Bh���w��TL��;���G�z���-�5h��#| ؿhSN`����")U-8y7��~GQ�n�x�$��8�u���#�R7�ش(�w༚�}(g�a��ꃵ8�� �5řt��yΠ'�;�	���!{�Ӵ g��&r4��T�Ƈ$�C$&��v1�����L*�$,���\�>��m�4�,���ε��U�b�ھ��`�Y�Xh�K��T A1nHa�JH�w��
c�F�|#L�s��QJ3B�KA�G�B��$�*W�8|OB^f��,c�����k4����&5�z�o� �	 <�9$�o�U��+q'�8�~���ک��V��a����;�I�l��0O�%'�6M�Lɮ#�ZN�E�\�d�i��ȟ��<�����,r�Ԛ��//^Î;uB����.	i��Ln�r`E�hC�G�bO����/-T�b�#�X��;&ْ�Z��y�_gC��$z~�aوu�%��J<�a߶�W�Q�Oޚ�Zҧ(6f�_�ÿ�x��&Rx/�̥/<>6�o��x�J���<��K.�ɽu]���kBn���2-�?�>���(	V����1PP��	O�A�݆���hIƏu���BS*���2
��VC��#�}+�ܵ�>����-������b��tq�sP\:�D	�m����o�I�PR)�j.����y+�Lv�WP#a������sG�kf�pi�u�7&�c?y���x�rKr���L`���dy�!X�#���'�n9C�t�����ʃw&��i\�F{(�	��^�U�M�oY�+E�IJ	��h�8m���͍�&��f��,����������}����Q�&�ݳKc���)t�>��§�{�m.;2k�B�������ܸs���}.-����#��к��Y�:�X��ᆕu �н ^Zjc������V=�_;�l׳��x�aXjw16|���e���xIJ��3/mY��b�Z�4�t�~*�Y f�*92e#�%��1�� �H�cm����k�J`�
�p�	��,�\�w����<`7�ߒ��1=R�v�B:(���g<Pm�wC��Sn��sN���G��(��bvjM+nS�	Sd|V}q���2�R�6q��\G��F��N�G]�ٴ#R�A����Ȁ�����r�K�ƙ�� ��w��tO��C�V*߼dJ�r����^1hI���b����"3��,�8�ɫN�\��Y�)v.��F�$��ν@}'�2�E$G5U�c��؆u�ѳ����������9�����-����?lDwo2\"�m(P]X��6���Xk#ј�;^���וD�K�A�-��y�N�V��QB����$D*13/��t]�!���@Țu�G�XCH9s@��	�E^$�1Qҷ�T�X�<�~���r���S���B���y�)\@���⤢���-�����ڔ�gU��I��r�u��\w�/��G�+B�Ϣ�����eG��
��t^����C}���}6�L�*Q��4R@�:m$*��-���1��h�cb�Nqf5��G�rџ64�����h}(",�_�9:š��S;	�+}���ɣ����]r�{t��v��Z��&�
���hُC��l��41���#g��O�����.w�p�0W�ۡV�4�Ѯ���Yb��Eo+c+"�~�&�j�
�;�XR�23�d��s�az)�܌m��V���ybį���#�����;���h��C
*i%K �#�Xɱ0��RP������ �HL=�d�J��R��bj�p����S^�6k��&ģ0���9�"��z[GL�rh���S�,^;�lJ�{��f��鋌�\�2�$k����f�I&p���U���r��<Z�D$��1�r��S�<��/���I2��Y���pF~����3lOG�*��,4/��le����.�
dp��y�Ŭ��]C8n�*7������e�"��"��yq��o�W�#] ��� ���ӌ�%���2H�`K8�[ԥ2$]�sϤ��j��X����Gl�B�IK�c�K���?�(O�N�~ca%��(e�"��y����)s�$y����d0
ť�$lc�a��	�#z�c݅]w�K�^Sϕ��F����Φhl �=@(�-76��5-���z��2SIC�QW�s�^���:��ǌ:w��)��4 ����<`
,�5��W�승��N)�@�=���Nm=íπ\ o��5_� ��� "xw�$N<�Sn^���Jh�����wק��US�@���4}�7A�J�4-Ǩ�O}�h���̤�P�$��2�����wy5IW����|��p$j)2ޛF��/!eXl���  Z�t�T"�5�������>�DH�,�dx�ѱI+/�a.ȣ�U�&:ɠ�e����Τ�Hͮ~�4��^'99�gz��W��W�ŧ��n%�d�֥��o*6�(*���=�8��Yo�m���_��}�'� I���ޟ��rޔ'$.�&x'�Rg��s��ġ3	�A*WtdƱ=!\���Ȅk.�^i���R�#Y�t�כE������Rk��Q���|;#��5u��W�y����J�-�Ϭ�os�ޞ������O���7���>CGzQ^_л�n�r��7Z?�|Q2op��-*��SG���K�~�ZldrD�R��?����4�g�Xb��;��p��V��H��yp���vK��zi�*^m�+�K�^{��/ۮ5K*�Ȕ�B d��-h��i��c
�J\�"��x8��͂����A�{N�(� S�tql8�G�-LU��4�Fk���/MN?��c����!h�1�j3ϕAHF`���0��s[u�ʝ�bE8��Jo��S��Д�K�i;��C�4�u[������S���/Vp��w�p$s�E�	��@���^-�𷄉lN�t�O��여�z��>� ��X4���N�\2}��tކ��re��y����J�*�@��G]O&����61&��>ݲ)S�����/���_="8�U&D�w�I���m)?m�]T�9�;���'�Ձ��l���j��鱊�E��A����uP�i@ނ<�zg5������zI�'�܁<�W��K.-V\�3��L�5�V��ϳQ��P~0��%G��B��!���+n���Ɋ�(��Y�z�1�听j.|��+\g`(��M�_!��J2�@ar&�-��]�VVJ�;5���-���x�1NmlgM��m�զ��L�����Q�.��~oh�1\9a�3JM�y��ߵ!�^
U��a���/§0-��:h<�å��f�hFhN�46Ů|�Fa�b�[()���×E��s�����.���B����!�$���@��PXW#̙p��@i�����l��?����zP��7���f��S���qU;�,Fq<?�R�4G�o�xi��i˓)��)����^<�T�5_"��è�{�!i�	DD��y�Dn��8�x0� �G���7_"��a���ː��`z��$��y4��p�"e��K.Y Z5���tY�1GL�r�0��v� �&t�:�ϡ�sςl�UN�$Y�����^g��nhXG�D����=�80�2�g���W)���-p��Ȟ�;3���@�n#�'�1~#�[�Gvȕ�N5�r?w�		Ԯ��e���,�e�H�y��"�is%=��1Q����,�N>��ΪQ�	�o�ԏ���3�_��ے�`�x��d�7�~��~�<�ܽ,�Ǉ���x�5n��#�mp��#��on*���ćX.��x`4uli`WbH�g��L/`��Mpߓ�O�N:��;�
�IJ@��ϕ�`)ur���GO-F1N�Wq�A��<FU��m*j�:�[{4w�t�����-cћoI���t5T�܎�8�B�՛G؟�Me!�󞩓R7�����j�����	d9En?UX+�1ؑ����u �8��Rv�v@B���4�����8f��8��`��Ƭo=�ȩ����p�F�i��SӯOXA���,�^Ɍm-hzF@a��/}-_�����P����J�Y։
�ϩ
Gil4��)r�Ֆ���w���]���He��JKb�Ŭ��D�6�KT�g|�tP��I�NϲȢC %HI%���r�9Wҋ��s"�I;��O�}���]<�&G�.�L�W�O�Cҥ%k�!S��o�����I�	�Kԁ|	�����H����eUQ����M�4�)�As��[q���Vs��G� b7c�?$�d��ڬ������G��SkQ��ҽ�v�����J ��s!����)�Z5�+���u
�=oG�,9��2�$`���IND{P�ݫv�C��C�VPOn9*⬴ͳX3�#Ad&v[�~,�-�`:ả�H{���~��~�d��J�o66)��k?c�����B��Sj!/�C/2%���>\,9��(��-�-�f:����c#�Hմ5D��>�,���=˦����8�Ü��L�� �mK|~�Yg�R�u*����p
��N��V�G�*�כ������u�	��J�Z$�ԍ���쯉U�{���1Bɀ<�lKz�x�N$V>��Qd������qK�:*ߢ+��`��ag���?�h�J�5)���RE7D
��e���ў�<�;�RּS}2�U��M��ˠ�6��ݜ�o�)�2n��ۏ���6Tkcz�,uE �朄��ޟ�GA�_��sc����Y�k���N�h�2l�0p	�T�v�Ϥ���	��\��H���9{��x{��� ��S[�,��:�ʿ h�GA�v��6K����,.s��G�Ŷ�t-�ܬ0�}��L�	����ߋj	�z���*8S��M� �՝��f�^�^q��=1�,�$�A�ߑy�'�@Ḍ��g���'�6���2ԫ����hG�M�(K��5B��!e�Rc_�(�т#�	��pQ��kR����a'�Zus6*Vbɼ#b��Cs5	��O�L�^k��EΪt�zctC�Bt.z��
�2L��vOAU�!���Z�q~pձ�MH���j�	6(�t�q�@�zN��&��)����)���̕��4}��>�)�k���`�v�i�U,����U�E��n��-!�@. �|�5ix�[>P�B����D��C��8[:mDe�p�ex �R0l���R�R�;��EC�|��M�9�~O��_���G��L�Li�/���K���?b<�~M�C(n_�͟����
��`��������<v����qhCÍ٩����ztL�	���G�t���-����?�T�Z�����Ikl�N�
;F%�M`����������#�QO�:{Kf�N��r�=���Ĭ�>W�7�FU�+��4�v��d�����3J�ҟs�׏k�����oi���\�����C7PeR.]UYF�v���)�(�M��$v}Mϳ�������.�t;�RH����I=gw|�æ�/3���Y�\�JOF���N\[��N������O�(q%<kɦ5>=�R5�ߩ�rG8�6f�[]h3vD��}��̶�mb
GqC1"��?��H������^T�����+�-����=�R>qQʠ��݂�3���Tg��W�p?�b�$�S�nN�iLTd!��戅���L�jln!nn�\+���;A$�a� �UX�~^�2�h8Ძ��&*%j,��9�y��HG�<��L������(�R��En�6�x��n�Ɠpe�K6��>6p�r�g�CJpm،;���Gv��(7Ań�I��&����(�/�W��Aڏ�H�\�S� �d��})�XkWS���,��Z^�E�n�荼:&Y����BԢ:����WO���-$��ЮE�<ku�&>H�C�>�mu��x�P���
���!��h���q�u�|8Ģm���?�8%�q=��+�|*�=y����y���8_����}�!��yƭ~�C��{��۫&׍qi��� �׽��0_G�b�9�P8 ��R����f�+�c���f-�t;�ii� �>�]D��Y̱�;�����Qs�l�6���}T�(�	�#aU��۪�&�oꟻ��>�ԃ6g��	>&�qsS��B��<�������CW�/�2e�3��ɎfJ�딷Q-�t