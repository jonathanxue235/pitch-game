��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V����hN=��a���)�硹<H��׮��`̼��D�g�;�mR�#rj��S��k@'�q�/�haQ��@ަ��m ����x�AB��9��ׁ4kDr�2�V����ល~�>E�4Yܨ'ۓW��<%�`�i��b��0�-l�Ggo#��2H-й�F��\<�m�]T� *Fg`m�H��3�����ԥ�Q�	#�}�����3��U��j���#�����}emkN�פ�G����kҎ�����]��ǵ��[������_p��(.4Ga��B���8��Y����Wr��p�0� �yE�o+b_q��LWw�[Cp�ĥ�
A�j��]$�����Neȋ���aB�5�'�RTZD�	S��AD�7�9]��Q�l"��w��� �����q�6�A���e�:�/���Sa����"j̥IS�X�xh	,��~�h'��9�%R
�--:û��%�����?�B��	x��T�Sk�,�aem��xu�>8Q
��?���Š[e.:�B����U0?M��Mf'k��6��0�y�7>4{e-u�"N)wM�Xg�&�j��!��/_h��ЇZ�N�������]�~qinӃj��syn����WP�����42-���iϢ��1�nXK_#+�%\��?�f����߽h$	5Q�::=��R"��ϢD����3�����h
����W�sHݩ)�[�&>�)Fyx�>�p���I�@q�]��*�_R�<[{���Z������������0w�h&�(����Ywh��h�5�p� ?��Q������`MG��+)#;f�};8�B���r�����튆<��](��T�X�������t�@`�ȡ9����	���߻���\q���,����q�ݕ$	.ôE � ����i�Lt����\���L�GV�ka�s#>{@�ؿ��oMාr�8�.ac�G�&�Oϗӷ�^��5�nM4��g��hQ!R�����smpAd54�ځ��%�_�xu����s�%®���p�m0�?� �ؖ�T���D�J��kv���?�v|��&#]�ַk?��,�ӛ��"��?�Ë��e �^��P�����?a1{���W�Y	$��F5ef˲�=�d�1
	P^��T�B�����V��a-=�:܂�?�0/Y�*--�-iT�N��}���לɗtLR�1�DLY��MI2�)����Iд�ϾX/��U��9�g�{��>��Z�h��E�V��~$���z��ة��I�G�j﫲�p~����0*��7��߆�3Js���Ԫ���v��z����H��e^�Y�+@SٷFn%�;�uu�u���I����qFϓ�4ҨD��"�.�D�P+�t�iz�p��6����?��߯�6�O�۳�ObOV��^h����t�SA}�_�\�W�1*��Ŗp���UO�����C�~S�K������2��-v�t�v��)6���y϶huq[�ᬎ�l�̓%/Oݼ#�ް-+V �	���3m:u��/���+6.M��ڟ���|k�K.�YU�pX���iٷr�a� ��a��`�O�&��k��x��]\`C�U�/k�����I���w���D}�*K�ɔ���u�ye��Y-pO��DX���ج��o P��,ˇ�H�Y���[�Vu���f�R$Z�fִ�0��D�ZT�a�F�p���+U�ϣ�}Wv=�N8s(I+��)I�Y ��_�V�V��	��ֲ$���խ }��F�>˷0�N7H
�]�8��X<cJ�1W-�M�E��k�F	+ c�F(o4�xc�mϤa���`�w�5��)���0z�[���q_��gR�l�u��5$�����ve���	6��Է{�(���j*�x�� ��t'cOtr�v���X�@�D�Sܳ|9��0�_�D؅W��?��C,`Z�.�������+-����Μ��Y{�ˉ) O=u@�ӝF�<��{�R�oh�w��n �zB���pĂ-�+"�n|�d�a��3���JV�X򖎓 R�����	�p�l����)�3UuЛ��~��4�H���ǘV�9�Ӯ��G@:	,<�[�
��0DR}�NI�u�SᘐDo7�ofY[�Z����߹#2�X \�0�U'��40ZMcs�.�B	��a �Z�;uĒk��h:,��.���3�1�0<�p�A;�E%G��FE�s�k	����~�}M4��M�6�Q��I�[aF�Q���!�z�0É�	ɾ���2��Z���qE��$Y��d�
�t��b̓����eO��`}��ղp:��	��Ǔ�F:/�g<�6r���0�v�vJ�w��I�c�G&z� |t�����,Yz`�΋�<���=�:�(2����L�u�e;���k�׾�<֪'�����+��E'{a
N9(C8��B�3������^�4����@kZ�<��bD�G�5|i��~CI��\g\`<d��b�f6L���&x��VJV����z����ێ�c'�,�H�Uj|���gN򨷲�#�����efK$�{}P�yBP{U	1)��J>��Z����
i�(V�5^�D�D�Gt>S�Eڂ^n��j6��a�EF���e�J��b)X��J0�/}���0b��m�A�҆�c�� �Nk�.�Oh�A��nH���l�:�P|:B|zZ1�۰�sQܐp?:\ ��p<0�P�� �<�,���H�O�(�}b�XY��`�/_�}U��{�ނÐ�"��md#�\��3��#�y8$hOog ͷ����$d�F����Tq��AHG$�T��M�Z&���S)IPI�(��hA��<h�;>����ڴ��a��V,��,����l����8����Q1(s,8�策N��K�8O����R�ra�T��h�X��0eh�Rf��'���<M��;�|���ڪF$�(�u��h�I�:��ҋ�šL�����&��(,5��L3��qa6I����w"c���{k��QqK�px��:���w?��SK�J��r�Gβ��n�J~i�0>�2;ε+c�P���[����p8��D ��\�L^B��e6�Ո�)��p�_+���N�'�^�'��.�#A1M�`%t�.S�
�%��~��r��SJ?���Mw{�vJ�w�˷��$h��;Ley�lP6�ʍ��+���j���_Qn�ѐt�S.��W?��?k�۳;��k�e���+_�6	�c2���������B�g����5�z�b|f�u�Fv��x�:լ)Ѭw��S4�.��qk�K�y�o4N���h}CO���mEeӳC���N���S��j�Y�:s�ߢ��v����a�T��d�h�sT��
])7��4�)ٌ�@���<�/~����,�u!٭� 5�k̅<��<��E;9�z���n�r��@��|�z��1�R�6��ⷍ$ۂ8(�V���0|��,!��(�������5W����)	�[l�-�(�.I�P�tbҌ�RA��t��j��ZK�.H�r�t�|�t�̢��2�f�B�{�iԇ��>����74[�3���vhH�q�D�����B�;o�Av�O}1w(�z<���KB$A1�񻴿�{����ʽIo�YW�w�'� C�W���I�����TѺ��݈�wIx�Dy��CV�<fX@	�>nk�L���H2`�h�·��j����un�g�����L��D.@�r3�8#b��tK'�%�*��Ms�h�~���t���"�ta�� �`�M����f5��ɱ�U�)&��^� ��~	ݬZx��[`[����0���,��$ ���c��������<~��L����اg��O�t��7 Iu��x�Xe�,�3߄_VFiCC�ղ�w��GV��Z�)���W���Q#d鵊����hi��p�������/g%��z-G�ڙ�3��{x�����9o�8u�XF�䭫�VWv6����Q�]����g�ѳǶ��d����@��o��}_M�F��Lɘ46�:ж@"�m�=�HK�Sy�o�{���u�"��#�3&=ξ*�=	O� l���]v/SCG��n��&�O	���%"����G�& ���-# ��P�h�"O�����o�}鼙N[�D��"mi֚Ũq����'A�N�%\!��9"y�dC=��X)�[��L�F,C�+15a<,�m?eM��#����׻���m�C���8Z�i�
}�CDR����$V�sU�X���G����T������mwh�ݳ�E���dp���K��/�y���3VxS��2d¹����_���R(��ԊA��X���7��S���e�A�<P��&���r��x8c�!FP�Л��|G(�A��?x���~�~�H��Q��'"S:ָ������)H�����ç�7��H~��Q�#�*Y��HZ�,p�B?.N�7*�!�ɜ�Y�R����8S��F-������4�&%!���A�N��L:�1P;0�����a~��s�~����W���^���G�W�O!!7\�������C�~e�S�Д=��D�؛��K��է�CO��&�P,G��()	�*'�@�3L�H3�%��ˡ�8�!�.%�
4�v�3�Kk����[.�A���[���>�Ly�1����?�?�x(��N�:a\��]��"�@Lʰ���|��}�慸m%"��ڳ_xq����m�+p�FH8Ќ��/�_{��ϳ=�We @<�G����)���0[D�W�2�wk����c����%�g��#p]��>�7��.�/�:5�JIU\b�ըFf��
o��)��t:C]�95��c�J��,�������ӝ��A���x�ϬR]�A��R�����h���y�{������4��2^
��n�r[���$�q�a��U�pG�*��*�m��|�5�A�3���ٰ�v�PSMo���3�0'�M|>���{�]IVm�/wuN��������W_�3&�);1^ȹ��uUPq�{'A�Vo~s�Ɇz)z����a�P�&��Oǰ��`���ۨ!4˙���;
,�ѷn��&�B:3㒪_m��ܫ?��뵲�$��T{�yq(gQ�^C��@{MN4��!�|���SK'�^��)ɐ����?��B,T?᫮%?���4}�mP��tJ*��
oGK��:R
�5�5e����P�M�h��#�J�@˳�ф�����6�R2�W2�3)nZq�(J��s`�z4Z?�0����X`�ϡE?T�J&��h��w'Fu�n�*ā��*mK�;GC����Z�,��;QO��ǅ�l��T�Gs=a=6(9�Ô�Aޯf�K�4}8��ϊ������9e����Aw
�Gl�?�D{#W�1]��Q�[b�<��
��[��<:�rz�¤t�#eFt�}pd�(ʽj�T��mj�*�\��.���.%2�V��Wi��osG�Wܯǿ���7�:�]F��|F۽��n4l���]N^~Ci���9����֪����n����z/0���We+	���V��<0�4�4X,�*��i-�&��u=X�s�2X��9���I�������1ƺ�����.�H�ac�	�n��@��S٧�'qf�yD��ȸE�}�gS��g\�O�3���ѣ]��F�eX]0��%����v�((�P���]��6w!��3`����!Z��$�./����x���L���r�!��;���_x� t�	������ϩ��B�3u����7��!���"�|ׅ���$�5��"�~�2ul5���(�(�Zڎ���4V|WV�cG ���Kj&���*{��l�su�ΰ@�p��O�k�j�7[�/����Z�`�!��VO��Q˻胳<�j�-�S}��[����4�F������=M�Á�&��^D�C���t��f6��fM�K� ;�c	<=M;�IE�W�f��*�����#x9�fc�����4��Vd�3�W�X��t�_��4�@�S�>ښ!�i�.�S'DMˡ�,�5[:���B�Nм�{_���p��J�)q�|���}*�|(��I*��b��tl�Oo}��Vؾ��2�W!�9�3Ũ�������X6F�e|����'�KK[�,��G˞�p�����㴱w���:�#v\5��]��d j�8�!�vms�Y��	�������3UEHU�פ{K��/����*�?�I��ޠ��|����F��yJ&�������U7[��f�㟗r�>u+�Ve���y_�?�A$%E�l�'��G@S��%�-��ۼ�j)��@�ߢTOB�MẮ(�À*k_<~?�*;3Θ��F�T�'��5���ث�d�|���֥F�.>�=&bv���
���B��m��ǫړ�<5��B�"�]��q��k�?X�CQ�[�G0�y���^�S�	V,��~I���h�����y��U:��6`�Ɗ���J��WD��]��*��%5�M@���KzN�X�:�4��f3H���dU|S]��2'2��c��P-w-��0f� ��X`%�EdVx�TDA)�,����Yw�����n��"^�Pu��jȉ���6�w�V2(�"g\��U��ۏ(�Z�4̇�:��&�2)�*�6C�Z�n#�V ��C�e����0���U�L�3{E}����J��oD5��Ä��y��NZ�a_���������!�Q�d�?�Ǭ���K;6�4�8j``���㷖"���S�WQ�M��U5c�|v���K��G�;��9���vU�MKr��e�Js(�~�ڎ�ڽ	���9	[ ;�1r{%XɣrU��OT���X]��X���h(z8�6��"�(�6��A%�^�ͳJ �@���n�>a
`���6����`�����j��Y��.�S�H�'R��D0W�]�3ٙ��d(�o?��a�$P`3�ZzlX�ϕ�9� �HQ)v�T�#���W�q��Dkp�C��:��\�:���=����|��r���A���Vr�4�-i?u�C�R7�C�Dt�>��{'k�ХwLscK���##k*����p�-�^Ф�U<.�`Q��S�����ӛ���e����iDER���d�2�f��(%�ټ=�YJ��Mxq�p(NWWס�ɗxž��Ͱ�熴�{1&��zɔ:��H�@���M��T�
?��ґ��B]w\�j�i�˭�UJ#EI8{z�Qn��W�TW
I���L~g3ѧ|� �u�_u!O�r���7�@B�x�����lwgB��#�o�K�o��߾@0������!u@q�J��٧Yy|R�^�6έ�2���Q�r?�%e	��X��c��'j4^?v�A�<�%�⟠�����6m�� �K%Yg�wzPl/�ԯn�pc19�X�1��!Z����)�������>�H���3cK�� Vp���D���~�6v.������Y����N�"4D�M:%c�B�c}+R6���7�����+*��	��З(������X���
�<�������B��~r���bT��}1cލ�vF$Ʌ�ƹ��j�)�ӳ"�^Jg}+Z�~N��@��$�t�U�H\N� F*���������YYӉ5[�������I�ۊ'G�\�~�M�y�
�~��-��Z����A\�	`.�19NAn���פ r��Sr�C��\X�s姾���ڲ}�x���G��p�nw�.���Go^r2 F���B߆�P+5��C��:�I`Ł�K�.�Z|_'dX�B�s5��.�z`��w���1�D���#bQ�>8sz�T�G�`�+_v��P0t�9|-5fհ���E&Yh�<]ըR�2����&L"1,��#�DK+�Ooܜh��7����aT�k�ƨ�ZB,"���J�S�)ivUݱN|����\�j�t���}�;��ms�a�wK�i�wcպ�-Z��0�%�М��c�*�}Y6�zBgʶ������3�F ޲R�7��^Wt�X{i��b�w�>hi�
�8[P���;#'��Yr��v'����Vr ;a��3fͽ���a�5��S�P���¬Di��ǂod��3�<��=���t�aq+
@�釤�]�:���������}h����n�g�p�o�>�dW'�6���#��_;�|��6>i!��u�]�	a��xLX�1n)+5Prϖګ�0P摳�g�:�PPp�N�;��4�Q����)����P�<"FNt>�JA�c��	%��)���+���h��L?D�}�NVUo�"�������$���ڙ -u;f2�Ui=u[s4����+��*��5s��F�/3�*=�9<G숌�iZ�A���U���&�FA��Ҡ�{���P��F�J�8.��C���T�^aYk��be]9[���UTuk��h�B�y��
O��_�^Gl0A�^I�0�s�7�{vl��2�.�z�|N7:5/*�	��|,���$BH���K�iK""kk�Ql}*��+l��; ?m��К�SEܗ�Di�6�DI6S���^V�E��2��o����?��?��[Mr���p�ì�m4�H)���;b�m"���d�Y|h];=���v�"�z��f�.����l������\�Yg�H�W:� (�e����l���[^����*M�k���X�[�^���&���(z(L�3����bGjut∮�?�
�uuD�c�҈�#�'w��3��YS)��=��u�I��&B�I�����r8Z7��߫q�:hg�F�����/#K{*��o�l���Q���=��:��ϵ�i��Wر�jZ1�" ��%�Z�zY�u[�S��zǖU%f���0��}0CBN�G��:�-��z;��ߒ�G5B馺<'  q��I^�l�����q+N��@J4����v�,];�n9F��rIBm00I�B�! Q������x�k{�����O�Oy��w9bޟiB�D(aװ�o�L��uM��"������F�0B.P�E������;�[L�aq����{k#�X������9�U�r���.f�D-�W&��6"'z��	�)B0[�0J�?��H�����Ep_Ÿbұk�w���#6e�K��F�JY�J3(�_t���j9br�l�8�pqB��#�l#��բ-F\��%������#���K~L����9�ԣ�Kǲ!�fC����'��9J�J��������9��U�����A�<fQ�R=��������&��y1�k�	�J��Y����L�����1����4:]L����C��Yh��E��G�s����^S4���E�m6C��p�/���;$�q���t��U ���U�m(�O��a��Ϫ�*��`*u���V��%�]�
H��&�
���<�ďr�� o�
��Xxy����|�c��ʩX�#��D��Bg��y�d�Rsv�7��z��FZ��EQᔲJ7u©����������Xߛ���p]��͍ċ�@7c����&$2pF�T��|ia�'h	U;��f��%�6�.H����A�.N��0� :1b�V�4�ˁ����V�ɀk"��Bf ���nE���Im��*����7��ۂ��*���hx^�+o8���H��is�}�%���(Z��s�i���յ|�|�F\v	?6�\��O����$l�,	��= lz���B��{�Z��� ��������G�׫�d7p&���4Zl������U��� Iu����A��賌�b��E�O!�=6��\ؓ��0|�n��6T
�!M� 9l ^�^�Z�5�����?����_7<�T�[)�;�#�>n.ਓ)d3��zk$l��y�Khe��V�z'z�A��;��*f�=�Ƕ�=S w��m����Yi��r,B-�����Y��ByU��Qr��p���{���E?2���a�[����r%bH��P�k�*�������HE�a�P�2�v\�J��B�'�����,٢Ѫ�)>��$�>f����,"fX��2��	�����2Ēn�jIq�%�U�8`R-5�A��
�3.܋j�N��{��5L�ՙ�#k�Ѥ�?�h%�r�N1��[����,0sJ�;u��)���kxB��K0���bg���Yxp��|>�LMϹ�jcvX��>�����&Z�X���[��Ny[�#�N�����&Qկ?�i�h93A�q4�ejcYc����9�Y��%8��h¾�]F�/�[�Ť�v�F(|�UgO����dge�H8��	J
���.�4d��� �I/��D�B�Hxݧ,�C���ZG����%���W�(���{�h��8��c}V�:bE�Q	�m��i�궈[̃S��'^�e3��h_������HCh�P���q�WMP�nZ�o���M��l��������W���v䴎$��K���"+�ɂ���[g';#���f5~��G�u ��<?6��lF!@0QrK����]�?WZ<D�D��2�˳�f�fG�&�����R���4_Ϻ�������J��K���İ��}3+��4��BR5(7<Q-�^�2��O���%�N��o�?H�����5�h@i��6�he���f�Xף��߹�Q�\��/9�����&�E(�0?%��PT&ДT���4�1.�:^.p�
����_�Y{��g�3YVcٛ:+ 2n5��%<�F��" ��%��:s��R�
�83̊�RĬ�I�B��U��J�e��f�MmR�tY��i���T�9��r�tI��edJ���f�:�g����۪b�Xu$a�\�]���B�(���C�C �)�r��q�7���Ym�?{��Y;���wx��찠������FT�	�}q�Uo5��ߐx"��3�6Z���wM?+y�c��
��13?��oԀ��­�D��w��Nk�C�����b�w�Q���њ�t	���Ԙ����L���Y�3�'~�pz,�PU$�E�ts�V��naT8�:�6�K�F���rD^w� ��l�����3[�(XO/��2�������O�ם�@ �>*����4x_��Ph�m�!U zfH��f/f/�^�&�r��|'�
5mˍ%"�ɢn�GBJ_� �n�	�U��53+#�}<M�$kA�T�ΊGRU����������ի� 
Ջ$.Vʀ){��KV5Hg��h��hg�}{=OP�֔�ޞDy0��FǑ��wxǥ^O�#e� 2;Uu�irc�Wƞer�nw�k���TM����2�d�`*Q�
����[=ap��PΒ�ղ~tj~���Ha�V!�%��j"K�Q̜��c���1I`d�Tf�-�!�?Ulb �,�2��c|�㹐�����߈�ɁJ梧�8���kS����h��ɹ�>�C�f��`�G�v��n�����-ُCU��sj
̪���;��]g�"d�~2}��C�����/D�آ�>���kC7T�-��|��]��)�> ��7��}y���F�'Ƅ�����5�9��{wH�S&r��C֍�����8b�"��+\�N�$A�u�))����[�5C:;k�����i�ƭ F ���|¡G�h�ET��|	cVm�2�|����^�<���hhOEGo��Wt�|��ٙ�kk�۰��l��Ѓ�dT�� ��x�L�E�O�:å��c�,M��:��V��{��ڰ�t)�Wd����[�#��_2~P���x��Fa���2h�lQ����b9㵡W��\�w�3�A\�k������#�b��TH�D�=��o�߲O:ΘD�u$� ��ˇ[���ܹ��	h���=�T�H@��x��M�/���d�SD����~��bc�x��_��lW�7m�.(�w=��c�*C{�I	��]|��B ��ǣ��?ܾ�6����C�ۘ/-CV"��]���@1���f�/u)-�	���u��4
�KS�^S����&u�F��m��
ȅ\~�
2=}y�����C���?�R-�j�ÃѦ�m@͒*�6D5��?ζ*�C����t�M�:T�iC5e�=,�@4����YB����yX�ւ�f�}��Q�a�]�^zu���y=�W+"]?�Ƴ[�	��oZb� k_�Y�h�r�*[}�����I P��t	m�A�(ƅ?�)�
���A���S�+��b����c�Q�=5̸�s�p	w(��[P��gg�H�<��Z��L�=��~��~c�s����z0�g�&�\[kh��x���
���S^-�2l�����bH�ܩ�`��������p��p'�:԰��-;����;�����uqI�w���E�q��Y*�ng%:H��!�w�Bs���Ʊ��1��?TE8�}�kN�jR�7�,����Ψ|6bf�Z?'���~���w�� ��*��{���a�W�YڐC��
"?h�D��J���ѹ'�uqYrDH8�3z��zitĴ��7���0��Um�i�Lz��ě�^>~�or�[�s�R��д|�i�ӫ)��
��Y�03��2���/)�N�2�öf�&� ����Mg�!������63y����jyG#l��	���s���^rވ����	<�&hN��3F������}6�?�<�n7�Y�р�E��,R���H}_)�_�-�]%P;2�ѢX��F����s�ϩ��L�#2�s�r��hU,e|�k�j�*.<�#�b�%���{���n;]GYtC���~�]Ny}��b����h���6�޽��kbi1'�,"!>f8�֨'�p\��`Ϝ�\Ĩ '�R�m	Pˎ���Nx*�>�#K�wJPW ��ϰ��XK���o%�|��w0C�=����L���r������95~�R��Ήn�=Ҽ�=1�v4�*�xw!DP�2IM�:0G~� d4�[���,s�7B#8�����=H�!}B���;!\4葴)il ���
��d,�����������}�%|{����=B5��5���3�o�־�L�ۿ���&�KB���LXڊ+��L�̠�3����5��
-@s-�_�}W�e�~�,��mbL�`l�ڶaJ<$M����D�^"�W�c�{^��=ǥ�|y;���]#�r�s�9~���~�b%LX�]��_U������7�xa���=[�7�����"�U�:��0z��e�<�Hf��� �~�
�z��f� ������ C��`��F#�iT�r�W�!�����lL�@�o�e�ۑ�.��LFe���˶�ƺ��?YV��~Ge���]8��9��Oi٠�A�ϙ��"ޑ�q� �d�����f���t��?�+�d蹼-"�	P��~D[����a��l9�F\�	�X���M������9i#��1�G��7u�����;.�\rr�{�e>P�TL#F����H~ڎ�i
��\�R1ku�-�L�=i�J�`	�{����ltG��)��Msѡt��go _�}�sw�o��kM�o�|�m����hu�m��@�\,�L�D��R��m�F[��ě�7G:���s�^A���yc��+ڋ�F���,Ȃo�VGD�t�K������=5�1�)��!W���6C g��"�d�YF#�LX|#��b�\��4���Hy��\�;1�	�DűĊ�_�u�vU�W���؜�����tOo����@Ԓ�_y�����y�l�	�S
}��AH�x�/=2	���]�m��C�zd���"�1�)��� ��_J�#u���M�5Ր�Y>/�����s<���j'`z{�w�!A����s@� ���� P�&^���Ek?#��u<�z��A��{+-�k� �mI�F���Ce@���D�N��B!��O�	2A��SyED�+���o�p�Q�-�$浖f�¹�}��p �ę�u�̿2K~�X�ƿ��}D�c�\��G�GYe�o|�����M�'�Ǆ�s��M^�x�9�$��W��P�:B��U��<n���i,G�F��fZܤ_�§�׿Q��Ma�%`p�&���<$���� ��,�0OE#O�I�9���r�
�/�kn�8)A&=;��_5^.j䘘ǻ��c\�&�>���;*3�S}���~KP
vֱ'�6�������H�a���T��ᗌ�SH,������IC�n�.FO���2��4 >�C�i,���ZSs�t�W8hW�"�~kv����a��ײ�~H
~ȧ5�R�s�ю�|�0:�e�+��s�\�/����7H'���s+3�h]�f��:?����B=�t@���zp�-��{'~���=ݗW5�i$�;��� s��sr��_� qBl"G�g�-��@�Z\|>>9���-�����>�z���T�*��C�;ѼlDs��_jJqy)���$u �>��u%�x�]j��X�	�x�p���e��ɒ	�#��s����(��s]���8+!��6y7rT���r��B���ω���S%J=�8?�E(�]�� �zx5���S���E���Z�<<�oZ[*��/�|�.X&�"^)�a��9��:>���M�5f�|�s���0�م���*e�һ��R[_Jn˦�(����
9�)�%#lv'�S�T��3.�ҾP��sC���Z��A=�ίo{����qD�Jm�_�E��	R|�Ԉ� \��J ��[3�"� ԅ�ܓ�i��H����^C�n�4e��բ�$P'�15�E��*hx���y�D�T��;�̪��Z=e�C~�A�Č�ȶ~��"�q�Qf#h���k�nӱ��'��6��~�3��,�\�r��U�~��[�.\�'���	��C��azLtRD�Ar�����^L�	}%����^�<�-?�\���}��<m����yS�ɀ���y���
�?X<���Kz�J��p�����,�������P�6�xܲ��I�i�L]k�XI�9��<m�-��$�Ke=�|ے!e�ؘ�-��Α�hDp�깎U�'�^�2�&�7���e��C/�j0d��o1��m;!C�W�~��Љ� }��AF+*T�WF�&5�̱�$�*�6Z�ˈ9�}�+�Σ����"��o�^LSJ�d���<dos��P�5�9@K�|��!|Q�����T��B�H����S���7P�|~%dt�/�r���e�l8�IrA>}�<�==!�Xoh#"��+9�pGn�'�����4U^�%[���{d��D֝�[ߊXP��MSN�m�$ �g�����ʽaF^�WV-~��N��m���BK�z�+�@�]/�U76)"+��-8�[P��֐n��\U�~]޴��$�=N����D�n�� ��_��j�Yzb}c�vw��{��H�#r`�;�����295��b�)����0�AWvZ���1A/*���WU��ԥ�|u�>>.g���2�����mz�.��~ϒTu��kk�Wr��2����GȌ��I�\�>{|��C�k_h9_ڰ��Oi_{�1b�Xeҷq�w�]�/58)�!����(��cl��Uk#���bC>��ǁ��_����({	[.Ήz�zi�_�b�&%L�����\�A���:�B���d$����H��R���?7�#�ƟBjC�[��4� @I	%���Y����*�h#n8ſp�������0�/,��$zƆ?������ZT�=�m����0�<�!|�w�v2�B^@���f{�M�'����
Qe���K�M:ͽ9B!
0��~��婦�O[�3���y�Q?<P�d����C��3O`�qR��`eK��T�,��S���_��	�{���?G)@���g�t��f��N�3�:o�qK�*$��"o'���5����^C ������v�i,������P�g�(@�Hg�F!�fʨ�cx��?�6��+�O�}`̹1Q��kͤ4_�Vy�5�5ŏ�!�6��J$���� �>G6�+�dM��?H(�␒���P�"H�N^��_/<�w��pIh���Ԧ��S)=HRO�w_�$��w��<0��g#YW�y��,����q�p%vG�S�	�����J!�}��	p��׋��W��zBKb+�},�:$���8=����t�揸4$S��+U���ګ
٥@g1Y�^�f�vȰi���t+H���*��T����2��,�Hn�xrw��c�j��;�)��������'O	M&����'u��h�r�[
����H<k%����_J~�T���ޤx�Y�B��2խ��T����]��֩��,(�N�B�X� �nr��_q��0;�ʕS� 2KI�)�x͌��J��{L�����?�s/,�w��o�ӻ���Z��[��$�ϊ�1�B�{������XJ�e��k;�@�����<��+H��r��0� ��1��^����W�\$�j*q��+�O-�M;Xpϗ���G����ھ�E7���zor���d��b���-��'��Qpv>��-�xF(�&���!�wq2C�7���s�ؽr꘹53T��T�^C��M��f���4�j��Δ��,�|Mo�b�ۯ��>����_������m��}�"�D�v#�~��.\�}O�9F����2Őq,y�l��z�ۋ�n�>#$KSMǇ���}�mF�`��n1�Ʌ�w�:��-J۝O�#p���w6��u�9Iy;l�C<E�4����U��P�i�:3yr^�(N�o��.���_5j�0�PH�&�������͝�I3��
�P�-�/�K��9��u�@�Bz���p�G� M��)�ǿo찭-:�U�I#V�M��
�θDQ�����O�g���Z�ʁ�M׎Z�(�Q��䬁��'&���g���-�Ш_~�	���]?�XCLԙ:-�5��r}��������"�s��U�GX,k�t��x��!��GU�I�����>.�����}M�%�;������J�^��l���>�J��zW7_�~?҃+�O�S1����Q�'�=U.�qr��ڮ� �J��3�Ni��Hq���SzC>�r�}�*x�q��m$%�eO�kH�+6�������+Q�@���ӟ�-PD��r��o��/��v)s)<i��SӨ|A��l�W隲�N���"w]'����
��.��[���d��ab[��zV]=�R�T��
��:���$P]�i���W2�Ý]���d�-�)F�3?�_oC�4��ޣ!s��զ�E�COu.�X��=���*�&mO݃C�?+#��Y`�v�͌C$���!�@�r4(3Y������?l4�~4������@�(/�,��]K��ny�3M��
m��d[74��-�E��u�ϙ�JJz�oNi�e�������O�"`x�*� ��S�i���q^P�R��;$�r9l�?�L4��|@z}���^�x�K��P�c�r�=2� 6�Б]~�����O���_\HF�B]�4t��N�R��9��% ⫸Jܞ4>�$�(},Qe#�X$(���W�=t�X�_��VN+םQ��q�W��L�Z1�l|_' ��I�^}^�p@\
=?يs}Ǆq(�G�����8j]g�'hUz���8��U���"�acP�(�UJ�is��B�&�5E4A�L�N"�֬��YD��"(Ɔ��^�]�ok�F)9u�4��|�Fk�,��C��Arg[��#'��lS��F�Q�ڛ�4 S�#@R,�z�~a4t�B����j֪�q�ѝ`�U��s�٬c�T�I���WP5�B�d#�>��Y�W������r"A�����cR*�����JY��\�l
0�~h�A�x e���WFl~�\0������+w�e��E��
ߚ���А�X��縎�N��2�9S�pN�܍|{c�5��i/pw��H��G��m��S�(�n�?h֎��;�	Z�H�M>���2�Wޞ�I�֥'qd�K���` �dن�.8�@��n2�h� 0#����:a�J{t2�0�"P�B{��Uz�d�N�G�ꗟqTĀ��.)6��� Wo������dhq����#���'E��Νw���bf^�t�0��M�UZ��/��t�w�<h���K��%i���A�Ш���7��Z���rs7��E��,3ē�h�r��9���0�`a�<SءKa3�v8��2F�?�6���=&'2��>M��u�9�xG���&C�_7��~�a�,����$qd�7#��b�@x���`��jX�p?)&Y����E9	�����f�r<��cʕ,�`���>i�m��5��Aa:������T�z�^`� }L(s���?�NJ�e���6�/���.̇��Z�naSq*�	�ξ������,?}G�I?]��W(R(���@|4Ƀ�,ӀqR��&� �wv��
R^���Y)/ʼ��&0x�t'ZJÔ%���q~��@��O�1MH�Kh����;�M�	�n�]�<�B��������'���/?��@�����6*�%�#�k��������^F�����ux�Q��g�u|��	x]\���Ja��E�������N�3�|�cGӺ-���Or:��	��?�+;V>�Γ���>�/_�
���D	�,7e�Sx*�α�c����r������*���"_�����TAu#��=��h���W����� �x��h�@�B�xVy�B�b�jK#�q�XU��k��~����V����u�-�z��?��%�O�u����/�pm��O �x���qN����x���P���۾�wb�*�]1����y�Ef��ki(��jOQA��R��ŉz�~6d�1�T>�dEk��11�?�뷎�E�4>�<�����b�Br��{}y������:p�����I[�|�+����O�5��u��m4��i�(���z�;H���T򢄆�4*?i�E�O��Q�X�N��]n���&�"2F��D5U�*�I�ɽ����������S}b~�ö���D�⸛�_�,a�s� ���qճ��O�(y���4���߯��8�����ʖ���<li��ug�*�\P�)2��N��i�N�j�eJ���p����Q�;>A��>tY"��:��E&��t�Mߜ#�t.hL��2�y�&�mb���14��" k�����dS����ES��8�)8��bZ�aR�v�%���g�<ʷ˩Q�!���X�l�/���d��{���o�J�}"e[��{n�ْ�y�[+�d�;���G���B8�e�:�=f�R��t�}3hA$�X���� >��-Nc3�������p1������Z���.�����U�+-�%N��(�a���#=t���.6ߨ{�|��Z�y�!:n�s0���`ڻ^yxV&zFF�&����'BБdm��UJso�=�����Q|��~��7�	X>n�4���'3�wҘ^-6��6�ͦ)�^�z# f
`�A^�޾s K�C���R�+���R!?��:z�B�I�q�2%?�<�Tƺ��]��"�����P��0,�3����/�-%�E�3�F��ۍ�I�5����D8�۷��'��<�mG���9���N��`���?*~6A��q9���T@j����ca�{��>�#�;�v�Hp���`L,���G�k�����W���^&��w��ײ�O�
�J��e���`]��/�eW�Π.u�D��"�R�?^uTۅ�@�i����]�8��7���c����*���gY6ث]/�ʒpɂ:LG�j8�`�9��6[��/9�1���$�`E��O�ڪ�A��d����r��ڍ��$�����ŀ2>��l�E ]�
fKW����T�+Z����غ��ro��"Մ8~��{u�Mrp��J��*s�b,%b��J��%�&r�8�S�k�@ȑ�m�ܨik�ң>f��ch>+�E�l�GK�|Ǎ���S�ݚ�c�1�P�����?����z��7�m�	L��<#��`�.N�qB"�<-����U6�(�i��AK�@��C�VI?a��7yVL7��\&�����b4<Ad�N`��t���O�Z��g֯�`@�2��">���N��/o����~��<)FT��k_�\'�-�d7�	�׶�b�j,a���L�B��.֗D�	QT�V���d��Zi�Q. >S���yM5j���Ѭ�ٵ�F��T���J#+��i*�;N(3�9�.�g��[Hg�K�i�c�'ڼi]%��Z��t`f�9�N�e�����W��v�6�7�;��L6!���hVXL��DE��^J40��9���%��sk8� �ޝ%��Z��N�o(���Q�'�$��`y9p�m��?`��sأ��p;d_V��.B������6�_5�*T(P�2,f5��ηpQ��J_Uџ'k��=��'�cڥ�P^U1��������j� �?j�g�Qg#J7٪�5��[A���_\9R�����)��%(U�֟�pF_!���9�e�gi���P�W�U
���"�H��D%��r�#jřL(�?���nQ����#0h|��<�f�q�5sz���J�v�����;���S6v�Z�J���)ߕ�zl
Z�)$�g�F���En��(�)�����j��<��D�ǭ��vN#��z��YvrQ���w�)�ǅ��yj�H��аbs���� �k�.��'�Sq���2�(d0ƁF�r�q��zʼ�����XI��4�A�+�G�����RV�*���ES��ɐ!-WԳ����,�L��0ц�G�V� �<��/X!±�sf����Ÿ�%N����K�8�v��7��Hy�f��0�n�Z��`�@�g�`����tbL?�jvu:f!k��iתY(�9���IR���z�y�=���ay�����n��(��r�^{��<s:��v����C��>��-�Lo���+�&o�H�:h0}�i2�4�t�Ko�r����݈��5�e����]�X�N��*ͣ�;�	&p��۝Тp�7�t��)>��+��	s��i�4V���$IH���*Ĝ�#������r��HR7&O��`ŒP_���^	�X�1���R��yS=�NR�7#�Vu4ո8����wտ��2�Q6��>z)4d�_5p.<��B�C���L������k�8���g�.��T�7d��Y�$��m#��M;�Ɗ��J�7�RUw �>,nT�Ύ�j�	b�n秸Z�L��&%�	�Slr� Z:�������V��rI�˿�ƄÔD=�T�_A�gH@�[��8�*�����o�?�c�u3��ʆ�iL�s[�4[�3kh��=�*��|;��@ˠm�a��T*��Ud���n�q,j)�%�GȻ%F:g}i7dj�SUI؅�r��ӧ��mͨ������F��"�0\� ���`?f]֏���]:�����L��?�� A�46�g ?���e �EXX��W"�k�YP���Tf�ryw#�u�@��bY����IJ�
T���t���l��V���^$��쪅BfW�?��b�e[g=��yVט�bB:dY�w�M(�~�>oʹ�v*C� ��{��E	g��ke����w	�hJ�ѥ�ٿ��TI���P�Бn�Ի��n��0J�E#��Ba "�pV؆*���aP�Ѝ�� �Eiۛ%��ŧ����̊ۼ������Fa[j��ѭo��-ˉ���c.�Q���R5'o\#�tH��f�J��������\�@� 	�� ���)�%;��K��|�R�8�2�\��Y��ϐ�B����l@|�M�@=���pa�=�ƛC˃���s��K^����;�{��=kNR�y�G�j`;������.��+^� PE�>���7��Mr��JSd�g�πqP�/Y�0	9���P�{�������0m��P��]&vj����^h�Z���;�'� Џ+����s��� ��������eo���F�M��後�����e��A�Pl�'�L(j���ڃf���`�Ë����K=Z[N��r���v?)o��*&����1x��9�5M��h�6�ֲ��z��C�=�3m8�	M�O�-?����'�O��󔱸�Xj�.�\�,�N�'L�G�}$�w�rY�ĸ̉膬8fel9�K�u������X�4-k�W�+<�̤cD�[u���.����J���L��N"m�����p׌���q���nb;&�W6�� �b�d+뎪����
��������
���ʮ�#!a� =ٖ��B|/N��CT���=�4��NJ�P����֭֋����J�ѐ1�iJ�%����^G}��XUm:@��dx��m�A�	9I�RU��_	�g'ݒ�Z�El���9Q�_v��J*>��kg�_#F�U�2݆x��6G���L�0�X��|J�׆� K-t��ro	�A�,�v$�D'4@!C/�"�8��6MR/��5:�]�h����L(��%��pX�)��u�Q�ھ&HG�������'I|�Tw3���3Ѻ٘:u8 	��m_�Ơ�%��W՜��vE��X)��3F�BUj;^Iӹez" ���(�zjq-^ ia�������}ܴE�l{�@��RN:�+$DX���0�p̽�:k��1��9�dh\�u��W� �}��1�T �E?��~�)[[�a`��?)pK>e(�d61$)�[��9j���B�T��y�k�k=��܂�!� y�}
/�籏^�s��� ��L��L�>�h5F P��({�:V�9"Z��/u�����G�D�}{����q]�q kZ�B��+�UN�|暅��pO�ѥ�ˇ��76��-n,w��RE��-��7�n�+[c���Қ�4S+���v�e���@Na~���ۏ,2J0�dYmD�X�t��>�_�'AAUfQ�����B���(��Q��9��<-JK<�qo���=�S��D9)b����èr_ ���S�q����$���YnI+U���'b�U���k�d�b$		Zr_"���	���4�j���m��?�ȩ��,����Һ���p.}�d�:_����ݸ�^�?�����u�J ���k�&-Ք�G��}{�x�x*��;up��������PɄ\:�H�YQ�z�9:�s��cB�[+  ci �Ҽ��f�:T�/�γV,�Y�s���̷��=2�oMc�m��7�=<���~ޝ6�i��G(]k�{�a������[L�]~�m�ٗ!C�݃?�j6J:9��,>b�Lur,*����x�I�=[4���	�T���� A����-\�(��d�	c��>��uS������4��̼�[���=�C&S�Ă"��"%�|hI�P�H����4tL�+D�ZF��_VpU���o���7 �"�o�;X�U:�~M�Y&�KqP�h�VJV��\����SQK�=@?O\-"`a5;_v�O��!��+f��Lu�#\f�Q���{�t�%��o��-��m���9����f���� ����\���Ӧ`����㳻�NC����2�s�z*�B>_���������מ5r�.aL#��wpD����_�O^�"�
h�����h�L<	tW��4:���M�z�a�%��DK����q�h��(�D&��9�Y�37k4����H�?�䯠�P����V���̴�>�8>G�X�BU���&������|	4�و#6�a$����>si��H����/q ��=�V/�\g0�<ە����+���]B��?p,��!Mb�XR.eCO�t��P�="�a�K�+�D��DR������{�@�jéɘ��k�Dz�iq>Ɖ��p����_T�i�SϚ����/µ7�+�n��tu���3�6W Q"��K_�~HH�ಞ����;]���P���@�����Y��缪��ʎ�0(�C7��0s������z�f�9n��Xhq��O)�Z3��*�?�8��)���K[#8�����	�a5��5?ԫ�
� ���^�%{.��i3�en���J֯eP6�q����N[����CՇ�bv(�B�;����%Ձ��}	b�6ç��X�,�#�*i6$nQhz�չӹ� v�:������C�����aM(2R���ōs�|@"�����=� TTXb$\kP��k�O�[ܚZ7g6�5����u��"g`��i��`y
�r%�/#t#q�	ثw& �X�פ��q�7S���U�k0�v.Ds�Vֿ�/R)�i=&��/��03P�����4UtF�6N�~��N~�MftA:�)�2je���9���t����A�0dPNof�/BkgfWe"�#�;g��h%]�L%>����
���i�2�R7W�V1;��ަ��Q��-����xH��m�`�����69�ߔ�\P{�%;N1�g3�"���0�&��VRR�X�����:�����̨�A`l@���;aM�>��V/,HϤ1��I��5�#ݿ$����O�R��e�"#Y��eS�b�0	5��D{	�n�U�ZU��w��ŕ8,y��!�UY� �,�J� ���184 B� ]����+8A}���� T'y��;��f4����ܟ�܉�+r�|6 �*��u����5�M��!"ԣ�*Nw�ɕ��Oݙ�"�|�0��Xu݌������^t53�����7p�E9�:�Ʃ��ʙ�B�Q�^~�5\�u������$2`�����"�}���ֲ�]?��[���v$m#D|j�9���	�L���N��<+���@�cN&�VOͷ����FP�.?^eB�<6ej�M��C%���)�<�����\ye	��@�Xq�Cq����18��^T �r�~JH�U"�)��]�C�EU5�UعEB�vQ2��=�����G����ņ�IU%N�)�����,5���\��a�L �b#���V��$��|�E�U~8�(8h͙�FV���$t׏^��e���0����tJnn�p(E���m]#�r���a��~ҩ)�U���z4�����4�Q���?'IS��$�Ģ{�C� 6|W�{[���?�5\.�lf��=��l�?�4 /�O��bK��LX�(wb��J�y�*0P�?��$oJZ��5~{�m�J�|��� �x�8Ɔ-��^#~+�&����z�����4�s>�]���e�_���+�=��WA
���Rz��!����ߣy����\xly�&��9d%r�G��׈q�,���D�F�,�1Ms��UU�s�ӶT%�M��/J�m�V��{����
�m�Y�g��5��J33�����Ї+-�L1,�áb��H1����_ػdX��a���2��Z?TH|-��/�ʟu/>�H�ZG#L�C��6�l���F;�h��o㘟 E��#*�$�͌ �A&����ē6���̳�U�:شp��A�Oi�����3C��C _�E�Z�Ǧ�=rđKfyѥ�O����Ƈ��;�~V����P�T�E��UR��k�6[|��R9臬f8�Z�i��&�p�$�Ll#>.�8�Iu�K�* ,���a��Á�6��]���v��_�n,��6Ư�j�%�g	�Ȁ��/����R�x��aO%�]+D�bf(�&��c�u���ln�I�_$�?(P.J�8R�{��$���}K/��/�ſ��|؈8�X~[Qj�֓��[_���/���Xů�Ui&�I���UC�Z����N��E�Y2��#[���I*3o�&ĵ�r�J���#ʳ�K����=�/{O;��X�xK��1ܵw��4��H�VM�@�v��6�SF�w��8�ۢWA����}��CHZ�.6�E[9v|VmU����o��"ɐX�-��i؜�@^J������v��@խ�Y�Q��t����<�@��_��%m�Zݎ,�鵬5'���'�)t��2[y�scl���F�N��<�n��UFR&�N�IX�����)j@����L�
U^�wH���`?���N:l%�?<%��R�6����G��Q��䶳�JY�C�w���Z�nfP��8��M�%��͓��&���^&b��J��!Ơʆ�ܶ�-��
�+���}���,mpq��|
�}5y���f땰	��R�`<�ǔO�(�zeT��ϱ�8�^ϰKkJ�4u��}FxG[�M�Q;(��ĠE��6�/T���wM�y��{| 6��sp���'��ʴ�f(�]1����\�Arp%��u`i���T�g�ɭ; ^�u�y�|���d�����Hͧ_'����c��Ej{i����~�����c3�-�ƅ����Yl3����W2�ʐč�Lc5��q�ѫ�vʕ?v38�Wl�=��U���1'�k���g�n�F��2n�-�����!_�b��E�ݠ.���?C��dJ[���b2��!_y3�gT;:_D5���5�/Ĕ��hr0�Ca�T�+�P����8��Sݧ3�J7j���oѤ��^�����V�i�TUb�����.�-�FV:����J���G�р�"|�P#�B�I�L��u��P{k�/�ﹰ8�#�������k'�3&T"#����_�`��_���3b�1N�Kgw0�D ����S�;��fK��ω���%���Ǳc�N1�F�G�ݶhy��0���@s�#��ϴu8$��*`��7QC@���5#J���
�-��q����ǙO��(��
�-��X!Ȱ�X2]�'tq��qj���p�}IH��k�Ae��z���p�^�mę2���Ŵ�X~��[r&Ic��@6��&�������b�����IR�����L�B��7���ː*�^����	)a�6	���;L:~�y!%�V��
��
�=*��/S�=�C(1`�N�ON�sqI����E&U��َ�m���nR�Td����B��c�5M�d����l�s�O���M����͙�J�2�<�{f͓�\8T�:�4W��G�b�M�3JW�����e���D�U�EQ7[��؄\���j� ���'��@�C�Do��[Jd����o2�Jҕ��>Q�)����i|4�z��B5����<�Ɲ!Qe�B�Z���=���}\y`MP�$�&3��7���ξK��5M�݉=B��X/�#+$z������2�R�I����a�'��
��tB�}����T<D�x��	�K���<�ܞ5���]���Y�Lv]zX���}�6CHKU��z� Q2FiJ���3xۑ�.�Q���Q�051ml���_9���v>|Gge���ޞ6[�ts�KaA^�ڰ�'-9�dX�S!���0U��9du�h���4ZJ|Kx��!�(�`e���B3�^��B�����"G]��Nۺ9�U�VBw+O���D52�e�����_P�`ԍ�#��'<D��e��y��nՂ!<iRK����5�	]Ti��$L��D�wp�Ӄ���D�+=`�]��pY{�Z��U���1�CӑvqQI��Z��|SP��Q��	yv��"3����,�;K�S8��E���lG��r@1�J�E%�&�dR��AbP��T�*���#�V��P����hc�J:�C�ŧ�D|/h'm�)�r� �Vt�� e����M[V��0���)��m�A���5W�(	iRn�S�Mf�y��-����jTc��p_�QK�(5ai$L�I�������t5�l�:�K�_zK}�<�xtϗ�-v�Q���������r{e"�ъ�͍߯d¸yɾ�x���+�5,+x'�sB��ø����߭���f�6���{	�� �`�/ׁ��v!)J�ҙK]}.&4��\E���)����H����\n���QG���*�I���w
@ h�����M�u�kC�PZ��9rW~�D�o�����ؗK�-�S�s��Ͼ���dn5�tU聰�d�(q���_W�?�"�ۿ���f��6"�N�����Z�Y������0^шn��[GI0٪R�uȯ�W�VS<_b9@��Z51.|�O#�b�8wG3:��(eY}!�XWeg�60�4Pu�`D�����������D�e7)}�7�ܵ�I������YlM:�H��`i��b�Grv�x�h�V�9�ʽ����6�ʘ.?nv�z_(���R&~-��.�v��$����:� AHr�f B��:�S�v��Zy�����9,.s���~���/��)էR�Q�]��q#�"�cT���\z�	 ����/�O������Q�2��i�K�f��k"���b@��Bj���4�<|п��~ ���v%Ԅ�P�.k5_1N����S�M*���~�/isf�#����0�v5ީA0'�������u"i��vە�1t��!^6�Y�3q	]�������c]�n�%��fX�����@E��q\��v�Q2\ �|C!�~ȣ��L�jQK�-%r����mNw�97���9��o�6�9V\�	�V����0�8�v�$�P�8��x�+�;�r���k��ՂBݵ ��۠z�b��9�Ά�`ݧ�1b �A�Z���f-��.F��>+ٌ�!��St�)U�Mr��*�1r�����pTP��৊���:��s�;�( �������3�����7ҭ�l��f����׶)���f�h2�0���/Ϥ���D]��}\��My{%��QV^gQ�����EE��Ή��`�Z-�X���?H�.}p�(_I�r��t*�wJ��ay��o^şFn��N��K%9@KTNeX�n���hyK����� g^����<�CW��&5'y=�����6�oST*�ST��1F��E��5�M ^(�Maꅈ��̨�vT�]��)_�T<��E&��I
��RMS�K!4��`k�C�@��w����/�r�R��F�YB;��@�_F�aCo�"�U�b�pxy�p U���=������pn�]����To�*�9Cfr>g
��7��m�m5"%Χc*�4A�Q,���R�qƀ��ƻW(�6߀Yd��	��N8Th��&{f8rn�Yp��@�|^+'��}j`�
z �^��Y6	F��z�N:]�]�&\s!�:��6���<+U����4�B�jlh���땥�æ�]�c�^�^�����]6A��:��Bx`c@�8����_���R�n�O3��F-=���$��3�?
�P�գ�0�Ve�<7,���w���eN#�)m�P�\�V��y����f���۰G�C2p0Zò�A���Ha;�z5�e�e]xUyNL����:!$��Έ���E�����3p��~?�B<Pco�kf�P�����\��N�[�[&�3�'�/%_��P���S��/��@���Yd����H���#%\���LԻ�E����؍�v���<���B�`M�PY�8`~�{�~�´<��"��|D��E�McO�t�I��a��ċ�>(�:ÌsxOMy:0����PE��*��7:�_Ґ��=���hgj��Q��;D�����e"�����{�����G�r�	�P2��jY���l))�6���=�K��a�d�א����K+�]Vk�^����w��Ҫ$���(9m��,�Z��Z7��X�[��m��r��	��;c�1��N�"r"H�G�)���"v�cȳ9�����j9T8j@~ɸ�3�.���2�h���n9
��.�D��(����ɢ�o�G~s5�4��*�('uT�h����9�R`p10g �Z���w��L�	U��gbI�Ķ�k���Q��K��+�2���%[�9�k��|��|=t-P�IK���TT����3�����>�N�"w�s�b�(=���oF��V�F�܍Nҩf�T�B��������.�ŰmL���O��8�1������	m}`J��S�UX�9x�7�V�.5P�筈[槉0����Q� �i+�Ke��A����
�퐈����f��^�nY�}F	�����f`�i�OjU���^���,`�초eJ�C#P�V	S���}D��鐦�ep��˵:V�����)�q��C��'���P�<=��h�\fb4t���ʄJ߰���%A���T�^���d\E��nu �ā��.y�'��nf�<Gp�����4R�?+=�f[ݑ,�Vn�?��Z?\JF�L����Ee�� 	�{$�b�z8�۬璇�G���x�wd{o�`�z�)�}t�Ok:D����՚�,�A=�ݨ �U��Fr�VFϴk�`�QS]��pB�3�SG�����_ NX�����p��74�^�i�}���0BŮ�Լ���g
���#y!�2��˟���S4^B-�PS�87:���sjH�Cd�D� �8�Jbq�U�z$3��ocp��?��#Z�I�S �aq:As7��7�"
'+��U ���V;��f�*�.��w�3I�JI'����Y)�?f��@r��2�Wm���(	j#�ώ`��ٕ}�.a�~Z��l�)��a����LA�/�Z����^.��d��z-u 3$mM��*}nh��J��G�T6E8{��[\���%>��N�^��r&��׀]�+�XP�Qki�>��Y����U;�a���9�eC{Pf����8(]/�w�_3�Т5D��S*�I����n����8U�Q�B;MDj��t����FD�{
�<"��A[촵E������Ok�|�����=� �)V3͉�B`r��{)X-�ǥA�!a�s�bxy��L ��z�O��b�����)�1/<x�'ny���ґYSm�T��N�� F��x�U(TM��#(x%͈1ȓE��/���f>����,ʷb��c��=A#d�H���B����k9������,4IK+����ѢS��aZ�b��t���Ki;S�`�k	,�E{jvCE����ȎTDo$"n��C�	'� ǾK��w�U�I�{ObX�]�%�!!�ρ�u�+|wa��*��4�^��Y\�����Mb�#�� "�#��CD�OǪ���?�1)�I��jh"��LrnCz4Oc��ܶ���rK�U��u*�G��w�u��1���,��&C�d�� ��+v��z��-�x�‍}�pl�G���.����1����AkpHnN1Q9k��{pF�(���GN�ݝ�YB��-3��<Q���j�����}7��سC�8�ҙ�o��`:\cG�K���Ń	!�(�а#1��`	���yg�?Dio�D%R&+Ŵ}�^F�Z2.��#A���|��A�+�N��)$��#�Y�W<���s��o���'�<��Hh���VʩChÞ7���(>f*R䏃����2i ���i�М�X8����.�3��k�}�t����D�s�)1TP����b>ī;c�NT��%�/&�Ƀ�h�sg��~���Ѐ�В��-�7�e]}
�������`|=��L�'wA�΄L��=pl��Kο=�|8Yl�����Ea�ޞa�G}�7�?y�ӄU���#��$F��ʳ������gOŸ����7�/yd�J��-&	2hL���W/}]�jH��%�Cv�>�S�x�����3-�
��`��8S)?�.��S�>��W̘�l{0S=*�K�\6qr����2�+X����Ys%�'
�=c�  |�6+��ŕ/n�TY!'��Z���,�ڋ̚#6�����x��S-��0@zz����W5�S�K�� ���4��_�p�T�Ɍ�o��ǡ<VQ���i�P�������v%�շ��R:7���� c���2>Y���wͬR׫?��:��d�����2�1���o�����$��S��irI�4؝�P���lE|��f�ʦ9r9}9z�����!�<~����e� �'*����� 0�k.Yw>���R#�Ӻ���iF���	@�4�T�vkx��^D���i��Nef��g��6��e���tw�A �YqB7l�Yl���RO�3v҆�T.�ؑ�-�%|���O��}��^�uC���{���U��{�����8���ˌ!����N��V{���׆\�z�t�:��x�^�X:��z3��r���r�2����=6��S����-j m:�I��#(�g�n�rR��)z8��S��e/&hG�j|����O�3C3��{�eK<F�1=z�}�]+`���`M=�ۋil��n�L{.oh�iO�Cr��
��-��+��b��O+K�e�캖�/l����@X=�۝ߩf���X� uq�h.f�k��ϯW�q*�KJ�I����[1�/�Ϙ�KX��wm�s?�+�%�m�霬���}���g�W��kC���te�J���)��
�%�Q��a�[�&�Sw�4D?�BW�vRz� �ad4�uiS�٢LM7�~&�b)�ǘ@zȾ��p;F����ʠ�gw�(�g%4�ʣ�پ�(�lxz�Cʿ��+�ê�c�9��5�����]��޻D�؅oP�$rj�l?5	q�H:g;�^6�H�T)���?�%�,u��;P"����xB������U����Q��w�W�/{��1k��0�j�݉]7�(#�>��QYd���<y����y�^^�	��66mW��멞@n���)������y�/I���iO��@�V2���x�y<�xvnR:v��H �Ɩ�u�n,R�8�4�hu %\#��o�� !�>�c��İ�iZ�?JE[8oxw*�|^�=(*�m=�:fN�uyA8O�9?|ur�?(�fE�3�n���fD�[��%�5*/��i�(]|�q�[5d/������b�9L�2�1��\ y.\�#��F�Tٓ㯾?x��\�\=�t�ٚ��g�9S��R�*���v���Z㼡�����76E�q/��*̆����A��/�A�>jQ�;��q�k_ǈ��TAeUS�vDlԐ�x�vB�C����³�	X�v/J�㴬��,5���1H���Y�n{��O����k�A��`Fl�Z��BĀS=�~2�4c/'��X"��Я�/���{��4���������eH�V:���l�ɱ|v�^>0L��۵L4��5���P͕vZ�O��B�,e�p\m^fy�x��LR�������Is-]�*��x�E�R�<c"�����e>1�x�x��Iҗ^i�׹&!d�G��՝��6c�n1�M�3R���q��6����H�t�,�!W=$,8ӯ������v�!9%��tM���Vq�lr�D�oĽ�Q�:�TZ>��z�&!.=��Dl؆�#����,���Q1??���*�++%z\y�B�w�S* �q�5���]uP�UV	�e�	�5V�>n�"���w��'�x���������"�=V�v��j9�)�~k4�i��@�����x��̚d�c<�ֻ�;����@)��	*�/M��1@N����&E�M}��w����FOb�V�=�i�!�'�������Ns���c����ėz٢3��-G�Ƽ�d�d��i�����q���<��]X�G��(�D��7���˽�ܣ+�0�M���q�׳u+�S�Û�d�iZ��+
_>���3���	L����g��@}fmE����;��_s^��{����U-�6��j�T�^>kΈ����� �wLI�E�ލ��x�i�V0���K[W��@[��2��hӖ�����ڽu9N���'!�4��R�A���X 0?^��5,�U�"�t��^e��7���<@]:�U�4����	��ֳZ�(�l�}"�T��]�㶖�?5u��<F��A��q!6)�"ק�$��ʎ����P�.��Ř�>�O��}�.%��y��A�V,{p�h������{��04#r�#��T)V�X�-��m1{ٝ�`�s�<�;$I�,�(��>Xg3�_�  ��c���A�J>6K�SeKB"ژ��*���-^R�E{�ɮ9�Î�]�|�yl� ��ڒW�zQ���a��ԍ����� ���FgE��B�$�z�x�ԴY���!��_�C��f�1�d+���tfD	b<3JݴRD(�.36}3ca(�>��E�o�jw�Y��~�Z'�x��>�0ZP�M��G���vz��eM�rwb�qm�_����<׈����FJ�wJ�sCu��k3�pl4n��,��Q�td�1��j7�-�i�&�.-��:R���^�uST]�?���F��FV����gԮ��k����&�_�W[8P+�������籧Fy����&U	���@T��S����-u�ħ��I�ǯX�	�~�z���OTz�~�֓` ��ؤ��P
I�j�N����0<>=bs�Yå�'�m�Ғ��}
�=+,61��a�������7}�wǱ�Eނ�J��v��J�Ꮔ�|,cã�����3��Va�zإ�ɤDI!`de[x �T1s ���F>�4��w��[	us����^-�\z=a�t�����,&C�Rp�|��_���ӝ��|A��i"{���`:�	Nx�v?K���5A2�*�Lv�K �'��tI¶�E��2��Mv{3'hK�꣹1�h�)g�:wQZN�C�����r�ی��+�wN���U^M�8� M�s�'�H����IC)�Y�P�0�Jx|����C�+�M���H��4�Y��C��cM�B�]d4����ҔH����g#�v�Т9ҟå��b�֠����}q9d�me���n_�̩��B�HK�j%�S�J뻁��'��X>�T���L��'�������гS �ݚ��	�Ph���9s��n3 cӽY+�v��h�j�H�`	��|3�QS�w����5�?w�ɩ�qxg��!�E��2�}��w��b[�����ep�����Zl��L�[Ī�	m�	�=Zpm,)9�Lq)<�oo'� ��S	H��9F2{4ᬦ��<���� �p$�t�%��4��/|4!z2C�	CNEbC^�1H�0'�kе��'���L�7�#�0��R��7��C�D��8�u3`��3����}�0���?q���蹷¹��L~0�SZHχ$s�CR-�q�F�ީ%���3%���E�uY��s�ך���'���ͮژy�/noC�)F&��BC�CꜪ��W�v�/Ԃ���lb����"���?�������pɸ�X�;�O�}	 �^���������+�|4��Q�����6��| �����xl�����F���o�n&����	b_���C�{�M$Y�6Foil�8\�|����zil4N���nI��x! 5I-�f:��W�<�k�����|�8��-�K����T�Wh���kށ��x��@�n&��DFS���\���ᖞ=����O��� �*C0�:'�q�y��Ә�$���h����|Ka��VQ�� L�Q#R���}��j�`��࿆ۘ1����}=��y��l�^ s�Q-�Po2V�1���\zn�Ob��ː�l��6T]hRLhW��v��x.w^��|OC����8\�N3%��]Dl1���G�W K�"s�v�TC�yJDU�b�$��X1��\M8?PU�G\zM��?X���N�T�k��i��b�i�����
7Xs��4�R�o��Sס_�`m)�m���V��㎼J92�~��`e��-�M���I)��s#f���Y\�2��cw=ٓ�(���:L),�i��ی�Q�}��J�.Mv�o��7�1�����@{�4��g�~�+Oz�W�./1�q���	�P�w)|j��R6 �%ӂ�G|B��o=�&�->�<dV�U�Q-��q!�ճAo;���Cc�����&��U�`�/�?c�#�<@=��cτ��pTg�?d�?e��y���"i���=YL$�
����ۋb��:Z3)!d�C�f��g+���q�鱁�`��u��B>���Ⴂ*�E�TL��d)����:B�K�Eu��zW��?D�G�˶^챿�'����i;bC3�yH�䃱GTwY��2*�NR�do���Z�&��$��ʜ�"F�k�iY������ճ$}�X������B���e4�z$�U6jϥ���[�c��%w�v���|��SX7�2Z���<ڗ
�=&�Ck#�#6f�#*�ȹ�
���4���{4j��Z�<gE�$�J$׃h�<QG��\nC ���:��ez7���J.����V��E�/Ic�/1B�m^�*,�X�cfQDv��cc�U�}������/4y��)R�������#���ln'v`��+�2U������"�F�	�=}ŉ�z��3�Oa�_���F{pX��zq�x�����Q�����y�\����W�Y	A�P� Ep��6a[Z�������ZŞ� .���`%�:�Q�V8=��Y�d�h�w^þ�kΒ�z���������� M�vO򕌵m�`絵����`���%R�z�(�E]��3˒J�sc���S�v�0�W�G�4��̘���_��dت�MX�q�
bbFX���x��Ǩ���L`Z�d3��C���EEm����L,�k����l���ΘjS�`f(���]=�΄ C����>��J�θ6�@O,l%���zش�8ʥ��5� ����o�l������._�U�]���>���ݗB��G�l�FS%�Z��o@��![:xv�ѽ㦋}8�!���B[�*,�J
�t]"�o�XZ�y�Xg6����{,�ֆe��C4��Ţ
]$�{����3��בU�b��M����I,���(g�*b4T:�H_��_Q��2����rg��±fp�6:l�-gʀB�Z������]��@��|� �R�/Ėٓ=B��YO����������YxA�)�^�'˼�QN36m�>2ĭ/��홼�1�VM$=���!k*��CYR��Ĥ��|(i���Y���?���bY[1,��f�sA2����H싪�NK4@d�� $=����͔ǅ�"��f�b|��5��:OLa��dTu���LE��)�SP?��E��
)��I��Gi�N+�O��;�_W@ڭM`��f�L7zCN\�:Z����l>W�m�V�-�|��@K�Ƈ��F�R\4��l�Wc��3�����>c!!�Qv��n��\�|��2�لG�S��
?�v/x=-��AfݼºD���F��Z/o}�Q���ַqI���g��i��j��qǟ���w�U���ӎlbZ����Z��x� V�=}���K�',��æHQ��Wf~r�W��G%�x�R!�KM�"#��r^�NA��E���2f��zϸ#6z��zYQ�`	f�5�`�'.=����7�����. � �m/�#v֊a�q@Aj��̓c�f��³J{k�yO���QQD��A4O�u��lx�+�C��9��K��<Ǒ������T	ύJQ�_�RuՇ�����'��+�p�P�v��9�Ι�N`����m����"���B��7qhDa�����o���2�P���lk1�e�-&�_?\q8D�ŗT���ʥ[�=Ǐ���[��73QRb�Kc�ȢR� *o��*Bi H8�c�P9������ȓ���8�V�9��P;�k�Y6��m2]�*��� *߄*o����ϙ� GlK�c7��U��..�I�ڗa�k*)�����:�/��&2�s�Z�E���Z�B?���ʨ����O��Xg�0mٹ0���<�"3�b��`����y�ՓOř�]?�ݫ��|��/~#��*��t�Ǎ5b6�h�!T�h2Oojc�2F�d<h�����K�#V[% W�/���EEd*�W'�WdJ>8]^@z���n(�X���'�ÎTPe���g�CϜ�I�R�g���f�-6���d<����	�؀�s�Y� ����^���L�em:�p� {���4�+j4�3}@��L���J}�yF�/���o�wт�E���A��������b�~62��$��*�g���iC<{a�UL��c�Z8���x�Ky�P�J�-�4��:�P�
�蛋ʖKbsc&���\!��_Byh��䎲I�.yn'-������Y�E���K]g��{��>tfI�%Oo���K&����ؘTP@����.����X�������$�u��@�f�=]�7�b�zo�p��a���d^�գ1��U$����� �:�w��v�a4����Gu7�"H���8��0?+2i���e
*z�M�:�P��\X�,U ���u߱�J>�G�x'�I�t2���l:��{�L������?�����f.q)!E�;���[n�BQkpjL�6��c���)pW�ܳ����������m@�a+4h���I�9*P��lM�DS�%.�v����:�&
�Y�ot<vD-�~"��X��YC��&��]�y�.k}�bQ��(����k-$a)�"�!�B::?�	�T�!�k�4��]P?�oM�Q[���l�U���0Y�DV}O}I������RX+�ֲl�l��6f��VF���X�aA��J�{�Am���Ĕ`���Q���QL�}՛+�Й��Պ���lm�R%�ƓM�l�)Nwc�I�.W�]���3��GXW��^H�~��{���N����-Ʀ�xݒ��Z����mɶ��$�����p;�fa��:Oa���M^�I��> ����s�q��)�V�ʃ�d5�ͽ$�Z���k���a,�*��ϝ/Ϙr�h��Ј���H����&�
+D�A;F���3�a&�ùsxn8�Ux�#X�'��&T�s�0��7�4Y'����-��|[�odFW��qt��K[�����A�6�n;��[P<��r 	����i�'�YX���2��5�
��+��}���f�u�ɤ�3h�;NzQU�w�<��O`Q>�g���p<$��+��ÊzgH�Wx c�c����C]�˳�F+����"�̳�iĐL��G0i�&�CGˬU�����u�2��"�VZ���W��?/Q-�`K��޹�f9�tLG���'V�Ŷ�<�!2�Д�ݗ�#��-���3+���*;	�-��"����gLy��x��1�f�x60�A��R����k`�����x��z7ᵾ6��M����a(���\&���S蚫F�9D���O��w� �pÎcm��p���`$����f���0q��2y����h���n3tɶB�G��*#�[O�<x�kRҪU�fcW����Xu���Φ��`�|�<�˖��+c)�������*�J�8�tP���)n�R_���*�jnk���I�P�83aM�.�IRZ�(gB�^�cC�H 
��q���,w�^	9y��3������~O���&P8�I�N��'���-i�K��[M3"֕hv�Y�LeU	�8ǡ3t]P�&�6}<�Kۿ1k-Æ]���x`~Jc/�~|����,1��S�V�����ӥv����M��]�k�Эk��V�ݎN5��ʹ�U�$q�LK"�]��	~�P6#�x��c8qA��=�H��v��U?��F�B�+A���Ŷ�߹z����͢~�?�o)Hǥz�&�Rv��8���ͤ�Um�`�Q%xyk/	Q��Wy�Y�-��K�U��%��H��-;7����1�JdwJ��Y?��
R%�ڡׄ#�]��>5�Rպ��@H���*��g��='�+c��"~r � ���.�m�q]�7��t�$+&h��L8�5����:�6��b�D7�.���W��x�U6�x���@)WvQMH8i���eQkI� H��Cx^�$�*�q$ܚA�Ɯ�W2�&�:Ɣ$�g9��\��./��g�Ár־���H��3ޯ�%���g-��62G�@L�^�/@�s���s>�0X���^^Dp�7������e�:ܑ�l��Z�N�?ʯ�X��9�FD69f��3ď�����?�w�f�Hs��X�h�H ���3��>H^4Ta�Ŀ��eEiV\�&�[�07tTB�9��nR��5�I�|��:��D�A��:�����sQ�t��z_��P++�\����+��9~21�g��O��1�w�µ��7���1eO�c�=T�v�2G,�'Cf�J˕O-�����xf.p|�����<���ǣ[C�቎j%��%?��Rm�<�f%|�/�J��4,�;����H���q �S��V�06��>a�4���0HyݰҞ�հ�b��,;j�ѫ6��R����u�Gs�u�~�0�0��}��ܻD�w��O��`7�yF���r��8���bhBߧ��XtN���x@H;֍�LS.q�?*������d>.P�uQ
�uHi�NK 'b��t��)���1���r��ZM_I/F5~PL_����_1��=tfUq�c�gP6�ߓ|�����#����o
� +���Gg���*x��B����Eem��	x6�ѡ���:EP�_�Ut7����J����#��_'���5Y�:��߄��8��t��g� ��z�X�k������3}������>��W�q�-�}hq�\�}-�2��ޫ����Z#����o**�S�,��^����W�K�Ί�B�&4�]�D)g�	V���s�8�O%�8p�����zjM�0)�f�����w@�J�f߯�eI���쟪/B��οv�ɉC���G�x��ɍ��O���(}��������(�mg/��g��8|�8�Y���YI�E�)��3!KQ]��I�U|X���t�>鯏��\�y�}<��u��V���:��i��WqN��&��D��4�f�.W`�n>OtϨ����#�����ʷGMJ��!"�W��a�p6\id���[�d�8m��?��y�N�2�$�RA ���SH�����(����
4���?Mfi�~"/@Rg,����l������:�l"��d�\�d�~�vc?t_G
~dot��vO��N�ԁ�<;���	� |$i�P����^�h����!1�(R�����[
T͟���z:�p����<C~���O{���ķ���Ȳ2� xf�E�}W"XbU�>�ǝ6kt����HX� ���.9����x�R�C |�b��u��g������&��$B@A���M,d�`X'$;������X�#�I�����$�0,�� g�#g\���>�upO�>mJ��}z�̱i�Y���@oL�$�y�6�I-u�ߐ�
  7��ƫ�[j��.�O�%B	O�g	y;޸��;VS>սnZ��+����L���~�̇7:c.e)d�m�u"�[�jf���㖋���5��K�g)���ɥ��ҭ�w&����aC#�^@t�r�r2�j�[�{=6�l��S{l���+:$dä[$n��z!�4j�Oe��>Q��AY}��5s+��.3�KB�$�����I�bYvh6�����!���v�cv���d�md֚q�X�k�W�����y�13�ٓ;mꅻ���"�ҥ54ށm���D��*���M���UWi���[Gk��ul����{�Y����I��!Y�m�<�4�T&�1�I����tq�w��T#�cݤ'D8�#��<�Ռ������1�����|��[������D1J���n뫌j�_lWg��b�I\����v�ң��~Ŭ�����^Q�w�*��-��F�l��\S���N����l����ɾ��W���~�oe����o�����?^�ŏ�U�N�S0�C�.v�����th�TU���,�AJ8�%qm։�������ǐ��./�yI�Pu$�!W!�G�v�Luh*TϘ_�e��4Z��
Z.�.~��<�n����E�\~�'���%���e�}dϵ�?.6J�>��F��� HdY3��Rn�Q�
�I�i{���,�"�3����R�flI��,�[HZM�ǝ����\̴/A�Cz��H{1�
C��泻�ȯjp�� 6�T����R�!v�����7B�ӏ��|�u����i�F�bC� "mJ�trP�ɉ.t+3�;���Gu�����>7M8�
�%`��ْ9�"��3��qF����u{�3�Ұد-�7;p�:�j@0q�Ǩ�r֔��k��s1Y���@�Ѓ�)��`
��b��N�x�֯'�^d�O�xM�c�/��
�q| x�e�(�y��	�yp�$�yx�N�M;ȋ�b�BH��0r2	��̲��AO��.�Kϕ���tF�!���`۬C<�,�hz��:ACr/L�h���d�꘱��0EQIt��r��6�Z��{�@v`�fcm��V�ˇw��b(u��R�����Ek`���	Fn[���Rt���h���tP] �m=���E���K��'�8�0&��NP5�A5��Ъ���"�c'�v�w�r~/�Ɗ����;pH��7�7�a����?5RS{��n���g#�!be�.K�Vۏg�m +�t��\q���e@��S�g����]"><RSl߶:j����dv<����;�	�"FB���_-$�7n�O��;w��npѽ���UT�� �G��R2����2,����Oᡎi'ٙ��(����Uð�v��>P�����S���>�j�ЧI,YV�&���;#�|rWC�^%c�.Qb���(n$K�k�%�v�(��Z�X�Y�a|c#��d]�8��>ߎ����)Kj��OP�`?#�Z"7����[Ȝ݂p�"u6�����b��O`���2�ÿ)�*Fq�-�ѷb�0��(\m?ێ<{�!g?\`�
�I^�]t�Ξ����JS���V��-�����1%��?� }��D$�H8�;4H��n�M#3Q�d"