module microphone (
    input logic clk,
    input logic reset,
    input logic [11:0] mic,

    output logic [9:0] mic_out
);

// TODO: Work on microphone 

assign mic_out = 250;

endmodule