��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V����hN=��a���)�硹<H��׮��`̼��D�g�;�mR�#rj��S��k@'�q�/�ha��pc�R�(��g�F�ו�����`d%D��G�qK�DW�+X���iv�O�O����9�t�0���`�<�F�2MGJ�g_Ю3����Na/��4-^}��ru1������>�9��& c�dN���(�lE#���f��; 2�{D�K��Ji���p��L�;������W��ˡ�M=\z�� d�<*ꖏ�<BP��g�,���r��o�֔A��*㏶M���$��#y�;�~�s��C�QDPfo�`��mʖ-���u�P�dRvf��V���%��A�5G��ap�Q�HjO��;�5���@�.�w���R�	"����&[a��A�=���l���LyBUN���<���7�#��KjuH̂�$�x��7	k�n���ӛew��9�ӞP_������g��Y�;�E����5e{#a�e���sd0}�������&�JpG.B��B������P#ϾV���>,�הAt��{�Ĳ�\��]�oІH�?۸Ӯ;r��+G}lP��-Ĝ�Ҡpp�h;i���iBl���;�掀��g>���,���� [Po���#9@EW��PW:&ovv��2��,4߃\Sz�=#EJ{�sχ�"1����w��Ō�.}V[�ۗ�!]��&�}���N����ݍƓ�'?���Ȓ�ܙhH�����_� -�A[[uuwgf�W׈�`������hf�v�ls�]e�;~��b��f����`v�K��

�G�3/��q���tY	���
_k��ZP�	�cգ�Ox7�cc��j?B������7�=��Qֵ]9�f�jy&���b�ѕ Q�:1�g���}�|o���_��*_��]^�{��fν���E��.����Q�{�W�:e�6]�j�:BR�E|�%ǳ�P�q� ˁ��Y���^Z��FQ���Ϗ�~�jt��	�Bc�rp�F,�����3����:�i�럃�p��h�U��XOU�Y=\1M���Z��L��n����q���d����;�}Ց�@��K��ʽP����$ݎdH�E�ɘG;�����#Z�jP2#A�sg23���be~b�m%�~���'S�d�M���{aF�.����ƈ��p��8��TtiZ-��䀀�n��H>�#��=��!	��O����S}�����(��!��҅#\�m����Ik˟�*s�f�\g,h0h��H�E%J�|#��r���b��:�!v�u�dv��ܼi�>c����~B0�]���@f	�E��hi����q�q��4��zb X�^cB�b�T� f�t�%�~��n�|j��	���3�R�P �
�Ћ�kϋ2|���gq�8��Z|�k��/���~&t��SX��%"�����tDNbK�r�?���1�w���v���Z?�K�ڈ��AU���Pc	0y�]U|�I���3T��='v`W�vh�8pkl\uz5X��,}Q�s��kL��s;FDĺ�޽��X���G6��N^F�$���٘�2��<���r�5tRc�*�1���ju1��]7�t�@$G��º��j�Y�c�+�kT�n�K_���Q��kUp��g�w��I���j�:�3v0�iɬSQ�<���E�,s�r⍉�xCE��f��T�e����0aS�@{W#�k��sE�TWbNY]f�߿�� M�1�@�8k����KJ�t(�TEDrt�n7�+|�9v�$�Y��I�k�z�����0h?�<K��'s	�|Ύ90��
�*��o�ʍ���QHt���.���,�dc(F���DF�A���d�}!H}j�a-����\C�c�[�E���1�]�������	��@p�.���,��اmFx0}<�'怯*Y��%���{�� �u$1��÷�.r���KS(c����afD���u��љ�=�0l�Nm�_I$J�IW�k�y� �udm���.�T�ː�!}��:-3�ˏq��A@ϻq,5�&�0?�!�-���|䱖,�9�v+0�(ɯ�ʱ,�Sm��E�<�aZ��f��&�B��+��W�'�Z��*�S�ǧ�ه�t������͢M	Ț}�u��F�-Œ�*7�����O�����½�lMM%����5�p6ꥭ^<ʡe`j`M� ���>��iƏ��$z@ZG���>H�F�k�Θ����

=z��5��|�T# �SQ/O�d0�Fc)qjg��_
.���M���������5��̙2e�v�&�Z*�\%k��]�C2�&��vJ�9)B�&i<-�͵�����^赵_��*�<���Qg��^X`�;�_��?��#u�ֳ���1�#4�ߊt�DR[�y��>�~�g�cF:�"Q���w|\�Y)��v��A�\��棻O+�QsW��Cȋ�)Kv�}
��8}�G�I�'���U��9B�ω[7^���p,x�N+i�j���դcgP��RY�2�kɚ���N'�Z����a���;���]k�E�8^�cd�+�J5Ϟ�[d�u8� �t$M)��L�^�x���e@Z+C�����_�r̲��D�<�!?M�+�����wY,�ůJ��zj�S��'�h�=�t��!�H�\%nH��D�$�
.r˴��-�b��=>��A�3O�]��_Rz�f!�c����BL����@�Qr�}z�f	��&�Л&o^�]u�|�rw�>#i!�}�ڣ7gd��9%o���������������Ƣi"�i������u���J~��Ƙ\�q��ҟ��2�tXF45��ک���IK�/�fe�[3�vo����uCя:�c��]�7.�5�k>k��s`a���L� ��WQ?*��Ӡ��T|�XLt*A馭����T��A���x��$י�iӝ5@A�;�e���E����̇_�-���w��V���cO�ƈRd���FJh�8¦-)p�eDX!��B��=�i��+�{���r��?�;ɐH�&	��W�g3�H���O?���vVW1��t	!R]^pS��Ĺ*f;q�9� �}�%~.V�gCⰐ�s�����Ӓ�����E�m�������" �`���qօ2���S�S����F3��1�"���k��fR귌`�i�O���3B�m��ݚ���+���*%Ɍoߪb;!�+��dW�[l�"h�ɻ�@�|��*y�}J�2���Aw��or���v��m�⛊���1�������0��&���(��1���@p����1�0�����
<�t��%��&�����co�e�F��R���Q����#��c�Ky��oi�8EXg��j,?q���%Y����sA��{5�)�\��|֔C�3�*m�n}N��?F��f��b��M�$%U`�-���9�
4�'r��|�4��<~ꮚ�gS#���1�@2Jm"��V�7��j�t��n7���E�
����.1��خ�<qN�HD�F��A�*CWo�PY�ݬ��G-���Z���L5^�V�A�&�����U��I3�T�g���־Y ���b���yq�,��=\���e����Z淕�����`�\�A}&���h5�Q�aK�,��`5(����=�@/|N�Ě��w�''
+�?��"����m�\����@�� ��>.	C�k�aX.q��є�~fv�,���uz{�K$FĘA�����;Ap~C�=2xi�Q�u�4��j����F�zOO��Mc�~��1Ϫ��	$�96�?ڞn�r�l�g���"��`y��6��>C��N<�B���z����ﱒ=�(i��0�|z`��i��N$9q��Z�k8���ێ�~տcC�S#� ��뮇�o��|e�Yf�ۈ>!+2� 4��1��MN����Q�y�};�`�|����,�� �*´�%uo�Y "�3�Q�I�Y^�_�̫A]�L�w1��1|D������@o��	�j��t�6M\=�`4e�����SZ4�A������
K��h!��~}ͩ�)�K��]S���mVf�����&��2y;�U����I�)B/��A)���h��Y�҉Toݟe�Eޙ�B�*�y�ٗQx�S�p �w��I�����<v�Ƞ^�˿R��>�)��/���%�'3 ��3�,)��T���͖:���8��C}oZ����ev��y�	�h*L��N�ľ1�b���	dX	�П�JK�9����-�h�
�<���C����یe�\���3!�7<C�Z�$�g�Wj�����w��h��'f&�<����W���tޯ�E���k������O��ڮ{�����������?�,~�ZC�����/��qF�]�%@��n
}~��*�r��� �i��g�
.׏�@fB��j�.q��4�g��!�H�Bl��o�szL	��3�4lc�X���p痒�b]T�R�'5�g��ʿtt��BHA�?�u䢣�(,S"�OB���;�{���o��t�Z�Ù��
�����3��窅�A0s̊��9��fR��3�F���yY�z�V�Ћ$�q��U����zb,���}�X�(%; ��=�~�Ȥ�H�<����tT��w(�\�[f��;�炢dvqM�W�<���\$�$'�.�qѸe��ݎľc]�^op��d4K��M���"��HxK0�D���?�u����j����[[ǀ��ҏM�ݫ.��(� )�6F���A���H�N���"�~!�J�đ��%�Kt�۴Q�*Y�N���nw>qJ�WA��&������Sab.�_�K�F'�mi��X'*f�n��썆[
�.�� ����@į��"$�^cJ��jZai�������\�i������,p5FUJ��H�O�e��g�,1�n��A��<����â��Ʃ�q��qS�bJ!k�MV���M�oXn�����	�<]�v�I�q��C��لv�
�
7Ns���2���H����h�f���������q�E?��Q�G;A�č����ߖ�'��]$#20��'���h��/���msǉ9���) ���2ۙ��z/ui���ic�?��,�Q�v���\����9p�\���#�LX�a��h#�N�E�N�'+����Ԃ��>���g�����M1�+�X�?*I�!agG�U��bK㕠�Uh�d)�ګ5���_K�.n!���{���%٨I�͏��)VOW��f�����C�M���������dy��š�S��%F� B[�����F����na�`�NL7��`�����?O�G���F���|�=�
�	�$A�����eX�<͡#�}���r���G)����R�n@�$]�.�%3k/��%[r;�͒fH����H� �
ށ�hU��)�u��i '�i�)�2�
�+��Q�qՎ�?r��LhB����