��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V����hN=��a���)�硹<H��׮��`̼��D�g�;�mR�#rj��S��k@'�q�/�ha��pc�R�(��g�F�ו�����`d%D��G�qK�DW�+X���iv�O�O����9�t�0���`�<�F�2MGJ�g_Ю3����Na/��4-^}��ru1������>�9��& c�dN���(�lE#�!��m��x����A�Ol�� ��;ˑ�<�A�+��}���R:0ʪ�7a���K^���j-������ؼQ*��k[�����RW�Ei�5N����T�0
}�z���E�v�a�_�� ��߮�72ګx��ysi7c��FA&�<V7Qf5&w���m��59�S�d��+f�YD�*/߯*�1�❨J\��ƣL0�_�ژS	��n�5\w����|��d�8v�3�F�-<L�����qLrp���7|y}�w����c~%�_-���1VMdKy��j��A��m��*���Q����e���g��?u ����G�N�e�e�A��#��^�z����+��X�m�����`zT�QT��}tA<�8�� 8o�Q^XݘrwGn:7�%;�}�ݼ�,Ȝ��@~D���3��o�1�9ߪY�����ݥ����tӷ4��o� Aš��'�8��L�1<�۶�O=��5���b��2�[��\�$���+ͮ�|8�3l��aa�l+�"|�[��mxdR80b�-�Pzy��9X����-oq���^����H��5p�����DЄ�m
�gB=�w�`�݇b���wSϕ\"$��q��E��>���lI=onÈ�Z��Ӥu4 eZr������皂U�����Э�]u���'G?����Y�;�q�Ի헖i<�I������=�*�T��G@�ЂdO�.yߡ�����J���+�!�MFN��b�ݝmN�f_����)Z�'0�1#�U�z_�Oky������B�rO+k,I�-4��M}��}�4)T.~F�V���56���X:��<�1��/��݆��R�Mp!���:�e�l�P�ʶ�EM��q�|�Fp���F~�d&�R�h}������� Lb�"�xR�.sK�i�h������=��]�
�����k�}Ģ�����)�.�PJI8����("nkO�Y��?9WV0�umVxo�CzH0�ڧ����y�Xn7��n`�����,4J�6��!$���}�?T�`���(����g?�@�����=�CN1 �~��<RU�d�ϸc�aP	��@=�B�s!���;��)���� �eGW���mXx�R�9�1�,�^������S1:��ma�Y���O�D����!hA�;Ɨ`�M�Q�^Q��W��׶��'�>�Zf�m�D�ʨTU"��v����6�w[�mH=v�N|��c�X�ۈ/Vh�c�/��[�k�C�ZLi��ࢗP��Q[A���yk2O��c���L!��=����:�괴ګ�*O��4>���K�ݕ���	Fz�{l������{�Rxb�Q*˭f��W;e*/ �F�!��H�a�{s6�}�ؿ�F8_IcE�۔�]K~<u��~D��-���]_h��ް���Te1��Q_<MI~���S{>*��N���9YH�Ļ�2S˫-�'������w��,Z���ga ���-s�\���N���~�Br��EX}�/c#t���hi����sѿ���Y�8 �5w=v�m��=fR<�m��mg�7�8�ذ�n̑)/u!GUN8z�[K�J�,hy�8\2I�M��'�Ixd�O��~��yǮ���륓Jˡ3ߺ뒤`1g
��.��f���/P:�J}w`F�>�NBP���W;��%Ƴśj���3�;O|c��|�	)���z��P8f1�I%�7�}U���d��.~��0�!z::{6J,*��G\.���@�X�w�Nܡ�\G�8Iz�/)��wK��&q���Z �	INġ��.'�(�|���T'��#E��i�Q��<�V����z埦��h�~�my�D"�����M@LPd~;����{^�
��$�ae�2�W���ptq�zˉ ��q�<m�S�Ԃ�x�� 8N?��[��)�� ��DhSN��+�Jm�0�����g֣A��{��pBp�O�Z^T��ˌ�e�?R֊f� <���֖�J�)~mVؙ�K<u�8�cv�*��X��s�h�8UK��F�s#�!�.�a&�S0a�-Qݓ��̢��PҲ�����$)����ח��?�h��^���naȎ��GoD��H�֋^���)�W9�^ u�׵��?�����"�X;
����B&@��N����B�ӑ(�s���f��|�r�y��Y�ʵ��!-#g:* �҂n���S~-�����^eޥ�����Nƀ�oR9w��Ui�HN�v�|pׁ۰�;�>l�s;�H��K0�M�f47�3m���8�Q�����k��Ǯ��;cÁ�"`E'VAи�3�:�������n���9�i��@�(�c��_���̑�报e%g�t4Z��7θ5{��R��Q(�,ۂ��)>��^��-����f��.�R���/ӒQo�5�TKV��^� WͲ�S�r�Ѩ�d�:=��t�XBae �7/L��Hc�-�;|3���
2s�(ÃJp��p�u�X��CSN��ݬ�T�-3�O!�a��T�W�d;�	���P���~��)a�?dg��	�?X��N�+������4�=����;~��<�v@2�3�<�4]������64�0�"���ג�:�NG���Oǻ��G�,�)�li"5ꃂa�Ƭ���a�`L��&:�/q]��ɬU��rvlv�R�.�V�/s�W��Hp�p��Q5_�Ԁ).#��W��4�N�(���G����3a�M�0W�_g1t��W��XD�Y����E�,�I�Ƞ�VR��ц!^��?�.�ԣ�DG�GO�-�@ܧ� �GP�e��cAP�ͥUĬj�Ӷ��7�]��u��j��9���d�#|8O`a���3�|fZ��P�{0�n:zf�� SQ�Jed�b�.0��U�{�{�����)4�f�F�R�����pGZ=�k��x�Ե�M���G�g+F	wtL��
��N���н)L��N)
Np��d$�+Q}sv��K���w�\��n�E�ag�j���*"�f�BPe(=mn
 t��-�J+�~c��Q��*��z�M�Z�Ɠ|�]�M�͊����9w<���]�� 2��*�'n��FI�y&���Q~�3]��9#��@m�S+rcz���;P�Wi�Q��<�3MF-fU8k(��"N<�1��7�us�3��?i,����^qK�	0:����f�:^>��6���m>�҄�i�;�NW�y���:�>{���[(��2�׿�s�ck�MZ����`I��"mŽ�x?&�q2�������F�*@�s�[�:NoS�F|fyl����7%�`��_���8B$K�*	� �œ�����G�j}�&~#_#�z九ɁB��6W�h��`O��NY�'��ρ���rdgUeFU7�z��c��I� ���a�R��"s��ŧS_]4� ��DJߎ�,E8'X#��W^7��|>���)��"V&��jP%8ѧ%�<���=x�-+��F۞�5�� �[I�ݓiWaa��
%"MKC[�mŵ{w�@vE�����0�N�|)�u	= C�����9�'�R�ǂ�׬\�L����e+|CID6�x�V�M���W;����ٗ�;yI�"���^穁�D��	��+3����ᗏ�ំxE0�請�v��$桷Nʒ�4E�u�ز�-���I=E���O��[�6��7�h�ZjY2�M��^��bJ��h��N79_6�U���,M�v���B@��)�z3o9���^r��͎������7��Ӫ�$��:�Pʬ%!�t|ex>��$y�;����O@N"��Jd�n�6):��n�W X�$F?P�?�qݰ��yÈ�0>���,S�;��kO.�� �j�R	�2�xӥ����E�7�ceږ�T�_9F�X��" �*e�#)�F[���Y�T���d��6���;�âd͏ �($$�|�i�A؀�KJ#Tѻ������֓�-<7�,k۫��H��:�.�
��cs�|`1��1b������k�e3�x�7�u�qVD��E�]4�����2{�6�����1�Qn��B�͍mH��+2b|��D�
Si:ko4S�Nw��zJ�[�\Ǥ��J�QTs�-��e�DX�W�*1�eo f��(�B��.�<���:p����J��9y-	ՉD�m+��P ���-���E������%����bX�����*A5�-V5h`o[`�X~Sv'�l�"Sz�r�	�p�Z.��N-(+��ֿ, 6��J=_���_#�#=|Ev�[�O�O��GT�n��,��LH�Y�N�.ó0�aF|�xT�T��|�@קi� V;�ɠ1(NA��1���lI9�&)M¥v�(��i�׍��o]�x�-����ѱo|驰[���:�O���I�@������(Hh���C4?ݦ>x/L�3���k�C�Z+�P��b-&�eU��q_.�`j�X�Kd0Y	R���u�;u��\��>��b��#"���F!�^^;쑾l1�u�"c�>.	^��dg�w2���] dOp��d<y� ����X��u�t�7��|�^���\�qB0�/�j����͹�[z[P�=혀s1,^��� p���,A���%N��p�=7:����ۏwZV�,�d�"�쯗zK�CTs�bE���ު!q�{�c�nVP�̊]�}�5�qH<�|ԋ�A4P���x�W9�'��0�q�z��7`BxF8W�!�j��R�\g]�s��V��g�v�bG��~�r�ѮW���Zw��*ԡd���AS��O���nJ��s����Rq�zp�z�2E:�%�u6���5c/U�=NƱ�W�M�	��{k>(����c�=Jd���a�(M=�&Zg��`�bo���i�-;f��a�T�'aJ�"���j����Q�/,�FW���
��< �z?�����d�Nw��[�f��{ �^H\�3���݄�ˈ:�rn�(V^�A�MFK�s����/8�&]��
0h�2g��r�G�S}5~Ir�ʪ9밥� �<�C�q,:�:ض5�A"��c�0	�,�?��>��%���^�������J�G�O>�-W���N�iQ�M���E{���Z�]p�?���u`ܺ�M�.�P��4�����n��`T�1CX�݅�"�r���L/E�SVE� ���C�w�~!���~I{�j��??�8���u:���Ge"b`��J���z�F�Om���"����o�a�y/�I�����gt�jB
MR��G5����}Z�5��`��<M����d�pLI�����և(�$�C����:�0�_�_���u"��4^-�=ӥ�GC��r۔ff��QtP��K;N�SE��{���$
�`�T�\A�)A��9���^VR�:����<�����ǒ�%D"JK��x���]�����#N�8�����LaY��S��(��+�d��Y?�!���Sؔ������73��=�������Uޮ�P���+�Հ-@���t�o��w����!��R���mK�u�!��-�ű��u�� ���u!	����~a��=C`]�Φ*�4�u��c=1�cq	� r8Zs�>TBR�Qw�'��̔f�AQ˝�� �ݨ���2-8�4�ƚ��ag@���m�hdw�'��#(;,���X��{_Y�yga&E��6�4��,HT�����@Q�S_�:�ۻ娣q̿�-a����T��Ï0��������!���Y�/ ��Ϛ�������!�cq̠��&�E�.�{3*d�^�/��է�[�U�r�K��I}��^�[|鍎��M��:d�S3W�ER�:]�J���F���>r���:.TAI���Q:�D��f��0
��38���%��
�e�+��1C�4�a+�b��u�N��p�#��/�[�>��Җh*>���v��)S=���kQ'\2�)T;��v�Xʦz2�����q�.F��vc�O�Q���t�t��N|ᾓc��I�s(��Q�X_*��4Ѷ�9�+����6������q�=���/�zT�rNQ�X���z]e<a�¾�@�>Ǚ�>ڼ#bm�aa�0��b�����$�:C�F�^>�l���U���x���Z��j�[C�8��{�}1�#�i�"%8�2K���D^[\�:���
��]\X��s�Gw�q�{�;
Vs%�K��B"{i�MH)A����ի�VL�lp��R\R����{ �ޕ;Uf��02g�%���m��d���.e�V<F&�3C^��b�q��J-�-��f�,s(z�8iF�b1��Ʊ�6�P7	��=�8����Cd�=���p��\������p.�4f�/Vy��>ǉ���d�[�^[�sz����ox�\�����{�c���/�ɍW�H}���$��f�W�; � ����z�=�d�U��捆j��J+�HˬZ-�8l�/�_F	�O��UR�ʙ~ɛ��)�V������ ԫE�4j���ֻ��v��b����;��
�}})d!-B�{��3�<��`+.�K;S�NvWM���w�򃊬��?�[���Ƹ�L޻�<h�DV��G	_��\s�dw�_:�e��.Zܣp���������W�I��w�����il4���>/('&M@��>!R�>�(4xvϻ$���.]��X��8��K3ڵ��3��I�����ۭmGi̛'σ������I��Ø���,��#[ژ0���)�w�N���Qs�&PzY0'
�T�i~�>:z�$���
��l���J^��LMC���/�2�[�|e��@��J��Lh���Q�䚀!9��(��O��V���*�D�lK����zF�%��o��IM�8k�!�osdw��`�H�r�UJ2�C�t۬��P�����m���D�����>b���4�GH��$����?C��.��	�!7��V߿NX�k3�@��ܚ��ߙ�@%�4��"�z����N���$0��g��Q��+��}x<}A�^ܑu���f�s`)�t������qD�h^�ʄ��dB-�vy"�"k��ʕg�"K�6f��D�R�ǁ��\N^�jV�DVvs9��tbzq�@۲7�z#b1��~Y�6ɓrb�a����J�AK��s���S�Ȫ	<�F#���5k�:X;�i�X�1�?�/�Q����L�̣��WI5	����< �x��"�щ�~�yFZY���2f��h�ݧV��ȁW��g�	����+v�X�@v�YA��F��,�A�t�֒
pA��]���K�a���{���E\.6�`_�Ԭl��=X�����NG���k��H�e���O�ʮN���������_����]4�yP3P�N�6`;�����6��� ��I	� ]�L�:�=w�F0���ڱ�1D�VV����>��9�>�B�0����)3��{��E�
�>�5�n�I�E�+v�B��j��Ăc���6��ڧ"�X���3��@��*"v�!+� n1Jӆ'?|�1���^�e�|��Z�2I��*��#+���Ъ�ɰD���4� u�����%� (�ҏ�=������KO�(��!��r�~G/��l��K��ҏWܞ�A�
8+������Ѵ�d��X�D�f�L`�J�>GG�-? ����Y>��#��Pw����z��=�l� ��HR�GSNzW��g�$S�C;DfI/se��"���$��kT���C,O7͌����E���9��-׸U3}xc��w(����ѽ���Ʃ��QF�^p��5��n0o�&�6��Iع�#���8&X'�	����*�8�I�nd_�`B��G��Bw
d D��rJ-�H�}�C��.�@�cI�d���Gd��`�D���цy�,_�J��Ԕ'���=�:aC��k1z���:�g^XD`���K>��kʘ1��Q�+Z��/�Lș�W�y{�s����3A�\�v�:@��2\x��t�>)��tDV��rR��3n��Ã���
�w&
n���c"&�=����Gs*q�ֱ�\�ȏ��X3�&QO���9~�"pC3K���G�0n� �sz0��'Ses�)O9� �-�'���O�.���@O^��qc4x��sb�;���//8��&� �"˲�+�m�
c��D�Xi�wD�f@�:zG@u֚����N�vZ�Y��/�
���j,�Rsu�y�	���wj����P<���k�g��]T�*�.���o$�4
3����>�K�7Pp5�k��'CăAK|�4��>[��`ML��hH���$n�e�� ���RV����+=2�����O�Ŀ��J;F� �����iT��d
�~H[p��r"ᘖ|
��tf�D�(�����Հ�d:��O8ad������y;���}��lz��y s�؛w�ɚ�C�,L�p���6��=�����ĸO>���vˉ�Me2�`1�M�'�k+ε6��M��N\ЋMȚ5˷';�>���/��B~��V���c>�}���Ψ?ש�T�E�g8��fA��ց�+2��Ք���D}����i
�H\؉�,���w�@��h""��K |�])W��=9��|X�ox�5� �%�'ע����v�6�R��u& �@�����/���3Jz۱�����+Q�%ao:��(,;j>D78��%$7�'h�ϴ�f��vJ����G�$���>�k��ѹ���Gʭ\]��c:<�E�:,.�6xQ؎�F�^��^�2�+&�U�K�S�y�Ne�U��1GAًJ���5߰��Rxj�Mq^���f��ì֓��宥U<ȫ`ُ�{�,�cc:Σ�N�{|��*e\����|iCFߴ���-���,`b�l8���\���c��o@IP����ì`�]E��{C�^�,��0w�䱬N�Rd�[4�k���ŕs*�;�{�� Oy��� `���w(��:l��֙bsdM1�
�^qe���>���{�O��8I�zz�����T&���0\�c8|��/����IcM�Z uzm�Xb���C��A�'_T�����1������I7�:Z�^�σ����aJ�CQ�E;zW�k��_����A��_��aK���4��`����a��_C��4�{����J�����p���+-@X.�[��H����Ӻ!}�@�ct����1M�[18��2�Q��.�E�8�,�����a���ޒ�__���`f���(��T��k4��	҄9-GU^�\R�-w3�o�.m��a<�:/*j����C9�t�X�	Eq������YA2Y�4o{��Β�PE�S�3EH�Q͵�z� �r�� O3�K����.��n�k��VZ~	�%���4��\��R��3n
a�Hgq7y��J��/���<�	B��[�4m��&xk��@l����<߈�2/�=h��"�8��2��yG���|�ø��s�OQM�[���j����hЖ%�L 7���i��D�K!y���{a�jna;�0�ݬ���]2�p�{��c�k;JX�HH�y�"�15M�E�5����^+��[���nz����J�%�#��i�T@j ��`�6ʞ�
b%x*�814�EX��E�@�/z6M���iˮ�����tm�9�a�4I��sh�ω���0���:�n�0�ţ�*)�bi��k���h�F�ߖ\��A�ؤ�1Z����V���Ȣ/1n.Y*�:�LA�L�p�['c��T3�P �Tk2+��]a�U�ۋ����m�ԟ�$��/�P��Aui.w-�SB�Q�����X�V��]�~��=Ǌ�%(�S^uC����l�$�W����#��o�m��ea!�ꮩ�x�nb�f�:�ֹ�� rh(�Ə�I�gc/A���3�f��OE�B*]j.k����V�㒪_!�5�H�
 1��ֹA7�:$s������>��e��C�ݸ��Jd�F���۸�ɠ�D�E^����/h�ƦDi;V��C���@'�A��y\�OE.D#=�ZFI||��5���7�%\��Ձ���(�0�A:ye�6fa��a�n���EW�����^���1"((�/���q� "�"1�a�IV�m�0t�1�[���ܾ���K�K����W�Pj�i��/rs�g:|Vw6�U	֝�\�2�hՐ�k�Q3�F7�!��1�������÷���t}}x�ֱ�M�ާ<q	[	�x�0;��BW���V��Ȣ%/�������|ݪR;����ºy�@扙�x<M=���A8�I���ݛv:����$3ΒdqO�O�=�'\Ȱ@l����aL3Q�3���e{xcw�8Y�$�V{�~-# �Y���ʧ�Nd�t���n���;7�m�p:���cCL�\��"TY`Ȫ>e�@�g�&�8�$?���1+�����E��+��BDh��6���5�\z��t�f���e�Ox��@������/~�3v�:_�"�m�e/8i�0���1�M1eQ7�=�}Q@y?}