��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V����hN=��a���)�硹<H��׮��`̼��D�g�;�mR�#rj��S��k@'�q�/�ha��pc�R�(��g�F�ו�����`d%D��G�qK�DW�+X���iv�O�O����9�t�0���`�<�F�2MGJ�g_Ю3����Na/��4-^}��ru1������>�9��& c�dN���(�lE#�)�<������8�1�,��0�#�(䂍q���%C���.O�q����t:�5�ֵ.�U�"ɼhH�̼�ȳ��d�D�mB��� #���Y�Y��j�%�ͼ����o�t ��t|c����=�4',?N"��I ���1��g��I{FթS���
~vaa�;�xZ%�";1� l���H�#,\xO��=��-� ����O��m�ǵ@�L��ɚ,�u��ʲ����F��껹�����Ff��ڒT��`W�԰�M.��� ���?�-����Nftot& �g�+k�`*�����N��`�OV�.��{��!��<�P����r9r�^���+�<ʔ����G;���x���q!e���$�B�>ՅQл����}���?��t◒V�P6��L�R��k6�ʼ�(O0I����s��}�x�n�᨝t���7R8��x�{ u�_Dņ
��|K�/�8�9�Qߟ�Z����0ދ�C'�����vJZO�Od���V~��
�G��Yj�k�iy����8O�"RF0ܩ�m��Pa�x�)���f�>]kV��{��^��ug>�a:`���My�s>��W�Z(P� ����������H3�f��u #?/�M�]KC������p����Oj+���,��E}y�f�ei5�)H�X�)�~ ��a��5	LF6a^��w��o��~�*OrHn8倐eK���+�:�N��A]0kt�{�Io������wϣd�K�~6��I'jP�R~�7�A�=K�8����7&������r�#���k���?n
�_�i�����0?��8��)[$�������Õ)�I�^����*r�����G��N ]����@6��pn��A_|��x�r�a�0�o��'D6���c���!�^hE��C���KW�����UB76;�z�R5�6��m!��ǃ̑�Ĝ`���b?s`g�*&�(xRX��:��'��G��F)�$�����fYЌW�,�N���%D�]�a~�=��&$� v��qk�\��"�L���ba�|,k�\��r/w� �I�Iu[\���c)��Rͤvk1�W�L������r�RG(;n�??^I�hڮNo[2A��Y��xԅ5�u�T�3n㺅�z�f��iNn%�爉��.ů��� �P/��+�[zASO՜;�!xs,�a� U���j	�a��1,�I��N%��vt�I7�J����
,֜�t�9��ޕ"��u�zg�!ý(yY�"��}�
Ě]�SD����%��#������L����G��:���qR^�؃�ד��H�"�~ơN��J\�E�WM{>1�g,�p�Fq+���Z;S,�C�9c9Sp�-�E1�gG[�r�s{��� #'K�5ml��uF��O�0F:r�N�j5ٍ_3����=�Ihp��%w�l�C����`�շ��'��Pg�U��5u/�C����_��A��z�s�
fu)t���e5�pS�vt��j^Ff6�E�G�8;4�Q,�9�c�Q&n-�b^�����iǔH�فҔ�\6l���kggb�n��_���V����)�w�՚˽W��j����f!�넹Y��q|���D�7
�ߞ�e�X�_$'�f���8���CՖA���8��p��f��Hq��X���WZq��|aËzφ&\`� �x���k�����L�ݸQ��p޹Ҏc����MvdKwA��ƽ�ō�f�c�^��yWo?��&�A�[��e	Z�H�&�P�i*��R�-H�9���\l-�^�b��sn�t����'é���cw�̊�l.8F
���HKy]D����h#��4M�{�a�����)����6~R�(� ��� xuq���\����O���b��A�(�w7]ٞb��%��q� GН�O�Ƞ�����[�"�*�K3���)2�3k��r�ɁyIS����@|����%��̽���w��xf���!y �<� �l��s���C����*�h�c]��h���5��7�������"��[�˃J���%��ݿm�v���uLF���̏��s��v�Tkk5r�&�{�������v��j���z�5-n��<���n�3�_l=�S6f*xA�?�|Ox�ůvUb� �H���)�!�$�Y��z	y�șھ�u%@xU��'����r�����mI{A��抦�l��e�P��Ĕ�� Ŋ�c\�[��z�^�[N��A�\�5���XA2d�(ss�~��Z��o�z 8%H0����ƌ���yu���όR��n��%P-��b��]*���B�gF��~�Z%�\Y�J�sf���f�l�+d�:Y�9rw�҉U���`�|[X��#�yґ����H--�p����I�1��WZ=iI�ci*�g+���Vo�>E�m4# WH�B�%>�t���	�!�h�-Ug�ML���Z3�rnm��\�8&U24����h�N1�F��e|�"ƧY�nh���Ɗ��)l}�#�D�s�Hf�f%mg�3߈nE���b�MWs�O�H]���˸� ��U��:���$ПWy߅5&&������~=����g:X��\ ������mY�Z�!ɿ���7MP�Z�ۯ��^:��V.\^�=Zo��
U��h����aZ��=UL����C��p�/u�Q�b����H�+]_�ej�WϽ`c�x��ch7��I:RYd�&vZ8��B����פ�H��C��f����J���[w�����T�%�Xᤖ]���|�j�K9��zW��P��6'*`��z��4#A����21E�"�6�@����D�T,�I� 9��J�N/va.�^[��&|,n�u8&q
����nz�K��?�Z�|�V��Ɛ$�!W�Iҭ��8�H7�B>�$�ъE_	o|rz�j�T-;��ドL+yM2���HoX=.eY���W\�Ӹ"�>��0��v��Ε�t���$�}�Fsw?7�Y��W�B��sz�˘f����zjF�Y,{n#�;�$�G�-��D��)$��d6ć�j��8�,5�VҴ�2nB���Z��*�x?)v"[\��Z���A����#EQ�7�]�ݶ#��\Z��>x8ǿ��򮫘�o��~�.�By)���]��(5��>Yb�?+����>,D�I�< N�*�B,������QkF�c��`��dr��r����f�_8��?���R�6��6Q͊�\�SquP��y�1�r���v���\6#գ1YN�ɽ=a����Ox^"�-���!v���/N��M��]�?ǣZ���G�s7S�$��P�z��l@?�z=���p9w$b���pNht����P���I��2�ѽo��]?G�4*I����L�D�\/4����5������(NX�a��^���������]ۮ�DW��W�4s�Y/_�U��&�oR��l�$�6WO}d�r�5�\�"��/�^��Ku�E��:��$�"�μ�F���q�?<9&pJH�8}j���6�;W(����`�$��	,�j7�#({ڽ�X�ӣ�z1&�T�`����%�<0%���'>Y�p.l}���J�ܳ^om�	|��Z�H&�����LX�~�E+<��2p-}d�=录&ڭ�"a��_ ����������yݰ^�]Aź��i��v�kd�/��iWb�C����Ai^S+���NE>.e(����A�4�dd8L��P�\�Υۆqg�q:��O�J	�����	�J�|&9NDi��Cg�ORPr����EC�m;� P��k;)TPU�	#a�#�s{OF{�۹�"��9�]ng�ެso��#�}ڍ�=8�d�k#Q��۲��4yl6���?�<_;,�W�<��qv�2vb��
R�}Z�5�/���	՚H47L������V�Eٖ�)"�it\ ����(��Q �y�l�k�w���r�/>������U�漮XeTJ���#�eأ�4D�h2��7��Mqs�c̐]r�LР;੻�9a.�{u�2+%��\���1�>nSu�j!����F�܆�HV�u�+(«Az���j�Ky�Ze�g!��4���A�I����v2l�LpM��x�))�n�3� ��k�����{v#R�ߺ���$���u���`b�&�����$��HQ&lo��od�c?gB�5e	���<݌�)�f�g��a𜞏b��B�}�� �@*]|S�X���]+D�[+���_s8Q�]�F�����]�t:��$D��(Ph���E�|!n��B��1&�J�nͳ���SI{˙���i��5�0E�5��b79��;A��o�A71A�ʤ��&{�LpO=�͢3�{U߼Z�%W�H�p0�@r2��)��9?�u�h�Ջg*'W&\l�}$��GB�!^�h�]=������,����0��8�I ��-�[*B��1����|�貖�����J�/&Bo�s�BmC�)���"�C���0�Cl������u�BZ�r�Kn9Ǒ2J�.J����̧$�r`M:hL�x�
\�ȴC�5�䃥L��z�ě�@3��d�?^v�i�<\�F���GlSO��)��"(P�?>ډÎ��Ig`�	MB!�ç���%OS�Ll��`�T 4AC�\�H`B��X�U�C)1�U.�V(�j�n��pa�Wb������#��'�i�p���YC������2{k��I��t4� E���d��T�|��)��6ņ���
Je��m����������a��bI�k�.>˼n|&uK�f`,Ǹ#���a6�� X��@���u4�8�� g���%+^������^f��'��2�(��?�ݑX�@ƾ�	��ݠ)���8���-��Y��WWe��q���i�>�%R}��!ezDv�/�D�M^��!Q�a�?4ؘQ�?	
��62i-n��w,����	�.ߞb�}\�t����IO�N"/.B�g�*=6)ʔtE
1AqmfL�벖j�KH�l����~Q��)rpm�Jy�9P�v��O��Q
~|�g�`%'�mm����z�z�"�'W�rW��|���aь!K���ŖA�`��;+��T��92�8��r-M�ȷÅ��������|0.�FШ6I�? ��\�:Ҽ!�N@�^�Ā/��[m�&�X	@�8s�i���;M���	���e����LT���.y�b���8�spn��</t-�ͱ�SUB�j]���#0'�AF0[F�@L��-���>\�Β�b���f��k�z��A�K��W8�����Ʊ��gﴐ��a����.O�@#REq�������2�2ʱ�Gy4C�$ ����=�:$��ؾ����!XbxF��)��$i���nj���֪qh-�����=vx�6���	�n�*
o��<�9P� 0�AM���s�R��<Ldϧp��ǖ���ay��I����Gk��_��}��,�����_P�a�@Ebғ�n�8�GCՑc��`K�I��#d�<�E�ҵ%���O`3����vj��쵨�㳡�W�ĕ0K����$��܋�o#�+E�l����Ls�ɿ�>"�'f������~�9�8�	0�o�*�E���i����]p	Mc��u���8%{�Btf^S�Br������%CZ �s��ݤjٮxo6�OC�Y)9�vIJgEJ��'9�@<q4�9ס]Bx�5j�}��P�2H� �M��7,��<�����}E sS�{W�L�EE���r�4�TǇ$��ް�c����"^��>�`��Q�㹹�ܳ�X�)v�eL���e1*+�oE�{b`�Oj��BV�%U:]1��~@OZ��hݦ��r��o8���Z��"�l����O$��4v�x��ߞ���pZ����d�Ws�c|���5��Z5����NA��w�l�����aX/~
��LCD7 "����Cb��u�Jc͟�1r !�4�*�����W��̨�3r@r���>�i�P�!�}r֖*�>��ஞ����2%r�ܓ��w#�g�^��,��p� NZ�SFSP�;��<��:�ހ:KN喇q��u�%fa�����]�w��]���mz����@��`Q�vE��)p��q[o�ZX�a����.��o��?tne`=3��{�v��2$���VguG~OЦ�K\V`��lO�%�p9+C~4cly{�����*L08I a��-��ۯ�����kG�$�¾{���;���Hv���x��Y�~L]9(�>��Ju�"��3��+>�Ԋ� ��ǻrhL(K�= T0q�s1�Y��+��`�p��Zx��>Y��${J�yS���f��w�`1��'5��Q�A���'�x3�3 2˙r �B��ʆ$��q""�� ��F��,KL�5e�I�"�P٤�9�mt��fO��yř�������j��d���*Z���Q�@�����3�t$�u#}��h�؀�.��ϼ��G*(GM��F���_9l@�iޑX���� �p\ A��R�� D����N�sja�ݓ��	@�����5w��k�����#͔�Db��J�3$�EXr��v&����&��L�1�����h��e"�2r����Oܷ4� 7R���`�������ޕG�Y�q��������l��/@����������^��5������{���^��
��a��3CjT��KR+Te�l[��7No����;%v	8��DPb�-3^�zCe��F�� ��?�&0�k��((G��jc;�F�,ȸU;�-@6���QP�]QC�8i2��m=��<�#\�8��p5X�xGa}�=FS5�P��Y���QG\�6;4{�بE�����e�;��ϭ�M��c�S6�K������5$�0f|��G�90Ф�x
-�V�6���Z@�L����6�p�!�
dtQ��'����r6��Gb���I	�ء� c�"���`Ro�����#�(���xgk�c�%�|i� �>�lVAq�B��t�+��
gƩ���[��iw�j�w�����F�7�C�):mK�+"�"��K̿�A<���d�MR�+{���7�z>�4d�Q��J���gE��wH��@B������3�w݄�7��ٖ�j��� 5b�k��(=�`&��r���� �7"��������TyL)�Cz�x���'�$x.��={ Dy?(ԧ𮵮�2�#q�� �8�x�im1����k������ꮶҚ���'�:{�J�HwQ����yk+�_F�a�&��ڗsن$��>������e�׿��ס�@ӝ�9���c�4�#���'�T�|�C`��"V+���s��	F�j(�6&u=sߨSI>-�瞘\`J��7f�Ӻ(e*�<*��E-�3t�aG����P�-_��K_	�\���n?�+.�ءR:���6e/� ��9�|﹮/=.��[�D��~s��'����wv�{1�$Q|jf;<�^
N(�R��_S�����/�����>�f�L"e��FQ�y�_��W��ϐ�^���0�\������g���;�<&����b�95\���Sr�1��-�����.٢����V>O%�[�g""�����9h��D�����F��.�ֵE�_�p������Ps�}7���QZ�R4�ΎD���v�afA~ w��v&��x��m��F�m��P��ف�D-w^�W?�k1y+^6�v���y���N��+���vg�i<6#����e[Ч��ȇ��czP�������228�e5�N��F=���z������(�ױZ�Wj��<�[�qc3���7����T�L��Rq\��q��.�8~r��tE>CV@բU����7�����K�"���������\!�٬���jA�h3W�QjHM��K�z�&�����@9�\�q徬}"=����YI���JU��Gl�.��gF�T�U�˫�5NX��B I��s�� z[��l���e��	Y���i�/E���T6�J
#�T="7Ȳ&k�4�>�*ՐuT��[�|����4'e䲛�v^�N��}Q����߽D5;�	�����?�>Ԥr������(�r��]�F���㮎�\�����2V�R��}�3��U�@�͢��:�ȑ�/�`_9>00J�j�� ��C�~�Wp6�.|M�B}��F�O����M��B����ǒS�R�h���޼�KՖ�=�J�!H=�S4�k�� ��$uL)A���:�(��$��	��	�}c̟�e�nɌ�x],s;\4�T�; (����5�r� 5�^�OwH~��{ᜭ�^�����!W�+*��`.lùx.��8 �hg4��Y:F���G��H-�v�;	ґ#P�K�鑾k�L�\.�E�����ɤwD7�4���5�7��$��bʥ��N5h�ad��C�=�{ywK,Lq{�Ag�H��j��R�j��/����ڔX��5�թt������Ò.T������HW�2�A1�3
]�?�Ԯ�r��i6�b�Pg�2��Pº�Z�RJ��e������Hb6��:s�Z���G��F�f[�*]ʹB��i���zQ�Ln��[�5�
��#Q]w��X� 3��5�<	��?sV'�����4ڸ6������tĘ�����}���'{fݤ�p#+'潒��i�����K�]�����!'�\����{�/>L�FA�u���"�=�C�V�a��߄cma�Jg��(�!jԊu#���s��\gz�ܬ��{���X�L��bV�H�x/�t6mHۙ�S7h��і\{>� ��j(�����RZ�P�7�?���%P���a��P��P�GF=�P9���1����hn�~#�V��D#���a�lG����h}�C�@�I�e���5#��Gl ����ʵ��YȈ7��VBahN��R��h� SP�)'���t�j~�M����+�S)!I��
�����w�(eD������}�a���G�4/��6�\+K@h���	���l���B=�	��K�&!�μ�	�2a�v�P�$W��I.H�zSO��Jy��8��ӣYQPX��" 5�i����+�{ͫ��I-2�7!��ƈ=���3Eϐ~NjBVx��~[ڻZ��%;��ٚ`9�E>6v��#N��������~-×�k�_L�0H�=�;�>#QZ0����KQ�  ��nn�NFA�=�.6s0��cpe�?	A���a�ʛ����:*�y�4��-/�����5�yTiNtO��[��Be{�S�n�.��� a�t���{6�Yj������KU��J�ՙ��,S"z��47U����쑕�
Y�y��}7��(y�}�Ws�t�JD��;Z��s�M�Ω��?[-u,9��`Ɩ���Ώ3��娆]L�Q&��ѹ�@&_�vy3�G�c<ݫa�|�|{Z� 0i. �V��':���_/��H�ʦ�޵��������WIG���ϴ	�{�m:mT�d�,N�R����?\��+J�Y�F�t�����= )�Y��-M��y�Z�F���7!��*��r�D����:�2�#>��	΋eIMfgʹy�l��A�����n��7n،��9�s��L�J�2 o��&>QҔ��8$I�j���z��|FPi��k3�w�!Ŀ|�O;�Q/I���qv��$��l�_`���17<��0�Xv���)�ܳbs�X3@ǃ��ŕT�&�w����� ��a�8i�U��R2mzBj8��y��j. �yb��_��\���Kʥ��l��B���>��sη/m�*4����*%\��]�`���� �k���p����F�0�Z,%+<�sqTq���(� U!��ҍ�|/b������w�`y%P<�>�N�vy!CV�L|=�&��G�6v�>�v�[2ԧ�`3e�I�q�ɋ~�ID,�B��J�V�@�Wm���s�����bEk�>�܉=pu��<H��6NYi9�E���M����=\�#ǖ����l�u�32$dPl% �%	�V�䁂9s�RX<���3Ъ�����g+���K����8	�x�7�	�z��X�F���C1	����1���t��N����>���Z�|�h�Vow��y޷Џj!���~>���ҭ�{��{E1�9Y�»��T�u�}C��W%��)��P�`{��g��8��x���y����� k`�mxsV&����2K��I�:>q����FfЃk��A�=�����h�w��x�"���5B�$أ�H�R���@U=a��m�T��C.2�0��*���eW�anݝD���{	F�Z���
�#ڕ9�CU�15D������ Y��:<��>s�5-�ց�J�B.B!�^�#m�PD3������_�Q��ȈL�\w$q�B1)4�+�.*�,�7}��"�f�n�<���a��^����|O��?�t0%���0�n��'���f��F��O��[�m�)��v��� x�%<�Q�~��P�>p�Nc��'�Z�F}�ʌ���*jS�|i�2#}W=9�-��"�j�b���<����}��[�b�Jr�IY���I8�ǔvWԖ��R"�*�_��~��,&��Ýl��)����>������7�6��ޏ<�;J��������t1.��Z��&O�x�KS�/�b�[7u��)r�n�xJ��uq܁t�ze�+̄}X���}hV��/��,��Lil:);8I�ܟT�I�8ջǭD1jo�3Ѝq�[��ſ�����Ǜ�2�m����}��z�D���.o0��:�z���{s��"�z.
�t	���y���l�,�i6W���c��gA��?�8�^�Kx�L�/|��Y�Tc�p*Ì���#m�p��\}��7
�hL��%
0���Z؄B�5�L]��b�U] ��!�%Rh������jC�qAٱ�}��>��|1����ts~J!��JonpS�2�V2���s'�фd���]������^/F0������
�f�ER5r}(l�S>T�φ@΃�[y�4��ok�����Y�te�W��_b/%�|�T1}V�1�ʸ��1O�"��vkˆ�����}*��hQא��T3�E��c��9���g��!*`_k~��cD:���T�f����5�dvȒS�=�=,<�����V��'��S�d4����9���b,0��r���,
T��`l
ď7r��GHڶ���;/���J^ˢ�S0e[��{[���<��XAq�Z��s�&��&{���������v>��*~(��x��*ni�	�"R��*�:��֎�M�s��?��p?O��7���8ϡq�a�w78���|{:A8�:�GC��7D�Uah�C̰Qz^�Ω<=�������%���h�UaO�y����RZ��@�L2s9�K��y���r,�&����;��˺���(��J1?�Wb��`�ҝ����6��
a@��D��$
6��y;'/�%������K��i�j/����Es�z�9���.\c�@;���\�sA��L.z�/�����ϯ�B(>g �Y�,6�����8Wzr5H{���h֮�@+�A�(�nh񏾬$��qHX/�Mu�6h���+�����ԗz�I5c�4x�W�]9&�gٌ��M]�nퟐy)귓R�2�h�=+ƻ����o���<%�M�)ܢ�x���<3�W��WV��l��^�BK��t��*ݔsD��8�HQ��ϐ����})J�F
뭊�tP!����JZ�llgiIO#~�H��h\��- ;�Ҫ�(ܾ TL��@�M��|��.�\��o4�W��]��[f�?����{���'�k
�H�A m�fC��Z��!�Uuɿ'P���؈a�E�7&kw�uTW���J�XP^�\R�B���+*�/S�� _h���nh,YF>�J���P`���DD�V��e3�Mؐg�Ea#)��51=|�^��I��py�OgE��GQµ�EpK�����:����.��{�����ve��e��]"v�1�L�����x�M���$�G�B*����'T�l��1�\K|.�-��N�&��.͟��a6f�^2�AM�h<5���,�K�Ѝ=��r�F��@�J7My`��]e�m9G2hh��'�J�c�lB	��C���A�=�����I�ʂ��e�0���uǅ8^��؝������[_R�:l?�K�������o�-0n�'���?��G�e)Sn?Jz�_-�5��"l��ph9��Aj�M�rU�$�߰:F�k���>�2~���Qusخ5^4�SkE���Wc��v&�<A,!+f�a���.m���Fv�$x88}�=>�T,��xטТ<e��l�M0�.�Vf�{x��F�d
�W첵���d�Z<OGіol�ĕ��w��$�W ��h��K j��vd]��eG���D��p-����aI6^����Q����v�B��+<���j��n��C������� AD������I`���㔃�.�=K��Ɗ�21�p	8�	�o�g��I�Mʹb	��voi�d}��i���U_Ub�&j\H3�ǟ�i�usY�$~ힴ����u�U�o�i�3wo�͛�������K����/?My�����A�~�����)��5�b&��qo��DSw�.�[M	��{B2��A����@i��kУb6m��Y)�C�C ���!�(��޵S}��@�l��нC/���[�f\��Q���P6:��0��� ��Pj��E�):PGy�1�ڙ����?����^�Fy�/���uQ�*ڍ��<G�y6��dYa�.	�7Y%>�T~d�T�m�}�d�;1�3~��˸�.��p�uT�|,��O��儬<�g�շ$�:�m0����ȳ��& �Nۆ����Q4w0[QK��s��O������ja�K�U���dd�5z����U���*7��:� }��|�� "�F��©����&��K�L���N��]���Vu}�?��H��sC(��if�*�P�j)"x!������a�=�֙4{0.]7~���Zu�=_�F��Mj��[��sdw̘Ċ ^ѻ]G#���}�Ƽ��mP�]?iO�c�	��	���������rIK6 �>}��ښ�BѠ�[i$	,�S��S�ؖ9<u�ؘ�Dn޶5�2�W\���| E{S.�0�A�S��^o���o^R��LH�����B�OR�O(�\[٢�}�?t�.G�����L�E���`��TW�m�U�z�f�Z�ލ���iPˁ�â���杧I���񊄚w̭m�u3E����6����E�g�����E�B����I�7��"��E 9�{� vA�$�CԮ�+�"���D+���"�ɥ��u������<Y�e;7a��T�˴x<�H�T�Q��z��w�a�'�x%E��*\Q��ѩ�9Oy�r�W7�	�!�a��lOg��t�etφ���4ۉ��ҹA���݀j�Qd�ѯ�@������a���0FC��Wg���muw�b���&�����5����՜͐��q`�G�۴�Nv�o%�ֺ�BEɺ��ԭ��"�-��?DfA�~W����t��)��ut{���2�)�ǖ��@Qe�)1���pXP߂DP���̓�&���x�-��6%fK$�:�Hu�@�[q]f;�-vl�x���@r�[�il�X��ٲ��[V9'�3�f�m�Vnz;�z�~-c����+sq���֖+@"iw%+ȗ_*�K%o�7�C!B>2 Mv�����g�K�՝7����8H�h�E�c
��e�j
�����������!�&~����s�L�l2J�ix�I'�`�I�]�N�vE��Μ�L�'X��v$��`�9��74�t B�VeP�3(�a��T��|���@2�hmD��;9�=�l��Y�v���()���/(�ت��4�g�)Z-W|�GM7S@g���a��#F��~��4L�0�h�W�3TC������*8W'�P�uY'b(�f�aϊ��ö��;
�� �zS IOt�B�*}��)H���F�?��P�)Vj��a�Z�3猽^��V��Aa��b��ʍ���������N���1d�*��m���*���+���hu0��`���U�:@��;����m;s�7xv��H�u�+S��6$�S}tV�3i��|�Mƚ�C�ᢀ����4���H}�}2�&�]�^��a��%��>n?��~k=VUZʇ����d�#��	;�:�	μ�n��HO H��'+.�ǝ����bǢ3�@�8�6�0Gf��|���kn�d^n)L�*�s��p�\yg��y���W�4i���(3���3� �����#�K��$��ƲT�'�ӷm�M)�2������i�|�^����k�����
�iT�.��g[� r��3�cq��ؼ���� ��״��8�2�.�Á���`�6sr��7���ʋ����|f�sm��E�M���u�>���uH��rz��;W�ُ��"�f"¥����1��Ȗ���֢��ceXS�����iw��Gxל�U<KO��)I���4���Lޣ��	B��{Ҋ�y�`y'񼑵r�F�SL͙��ZV,�����(c�����|�W]�]dM ��*�R��9���zk`�)S�f���l]>�z���e{��n��� [�Q���G<`c�%#��?��ù/.w&�\X(~�%��8��
���WO'�jM��C�Q�9�������z䴾T� �N��vM��U��v��1_�ɥ��T�Ec���}��X`��j�"�����M�Z��Jdo5@����ӵE�.����6����b�@���'�63�M�(�nd��u�8�F��k�;���]u�W�8~\-��Q�lu�����Ms��jt�>	,k �3�ȉl�B����0������P��2Jd�{���:�U	��؛�, ͬ��1˶F�d'?߆�#>f���HC<oN]7qF屃�T��eOh����K�A�h
�����F!'f����]Q�&��C�"��ԯ��%{�a��S4�3���i�0#HU3��;��FոrAy+\kykb]����<J�^�O�#*:�%'[m`wNjܙ$"o��pɆ��s��9j�c>~g����X;��XҼ���֎�#��,�������)tdm6{���O�?㺯��UUC�����K���C��M�"8������>!��*�9K���h��
���;��� �v�*��h��Z؞���"�5��X�@-�����{_����O���K��}�����8�w������xR��`�-� ����;�0���e-	H���|$񊜥ANX�3�t�pË�42Mf��;�f��?�B���ORi�=�X�&�`!?Z@=�o)��n��㳭0��*�+t�3v�����7�1B�M�8?�/��nn����O=�GUuDK�.wNE��2��%�O{����I	{ɡ7�x��8Z�L�]k��\R%M��Ba��:��Q��l�L�C�~����m�'��vScۚ�Pm�#�Q�;V��̀c*�drR�NB����}sݴ^K�͚9iW2�������,���	<�6k���O���Ɣ=q���;���W�"^XA��.dhnٖ�`�JK�Ey�K����X`[��׊��[G�}�e�?��%�+Qh�	k@�Ȁ*���FUex��c�v]��!��x��Ӛ^G+��|Op��f�v�:fM�t�;��5�H�g�)/0��V��iBE2Q's�� �C~Qm���@kƚ�
~1`R��6�&$;��ɘ���;]�?��-�w�u�Q��Ҫ�D�̴L�K)���Dl��q{�p��gŷ�ۛQ�>p�ߦx_�B�z��&�G������/���Ҡ�Hl�\��9Pl��2��1����Gk�Ґ ��F��̴�8Ă��j���f.oŦJ@�D���aG���Drw�W������������Y�n]��Q%��@��3g2 �w3b-eO3��]<�����PWp�c�����w��-��b��@�@���[!8d~̚#�#㷖ΟФ �� �m�������D�X�i��A͢�K���/$@! Gy��Y����B��;8a�W�â�T��1n/��{I[����C��V�Z�ҔbuYI~�k�=q����;	�Qu(�8-����}z�����*��!�#�����u�B�M��Ѫ�y7��Y{<��6�<�9E)$����z�?�	�k*x�@�q�(�&�q\C�^���pu�5o������M��]��� un	� !�Ap�M�-�������IS�<�Z˄����c,�=����6���t3���?9X�ւ���ʢ�\hV,5f��_�����TIt���D�_ki2t;��U04^��0y���0�kml��	X'0�Y	�Մ���h�|[���u�j^�����fH��_?C�s�N�	���v�^�f�����KД������#�D@-���n襕?���rrf;K2�I�|�kN�m�C���GD{n����,V�>?�2�9����5p׮�/|׫���&q��{A�����}p�7�����eV���5@�W���������!����E;Q ^�(,�Ϲ٨��=�Ѡ�	��pη��2�cNΓ<���G���(bɸV� 1��b[���L�
�%�5O��-�r�,�O�8vWXJ7� �) �
�l���,.����*��$�b!^h���PF���:�BM�]���M>�W�zb��@k=m�>-���|�eCR����p,��ex�i�$!o���xM�_���^�������1"�OW&й��1`�Z������y>����)v��)5K��>�
���y���a��y��X�+�k%�R���y�Q?I��4G��������tU�v����-�;�T�U%�!o�W��Uu�5ܰP5I_��D1B��\
y,��}Y!�)��|7N�/]�M� ��f���k�)������C��+�Ǖ�����br�E7G�QNE+�IPi��"� �[t�L"{2�����ƒ��7��O�¥'�qvIXϖ����>�b�B������Rq��hu�)�����]�������=���-�(�R�29"0������b+�X�XR�n�J���4tT�s�>c�pf��J�r�G<����BTYݣ�{|@�&�Y���%��e�b�q�WgWэ4���`r��n͜�u����<!�?�.e��r����	�0�ڔ���-�^�~�ҽ��u=�[�S��=���	�G�<	\�V?}�#T7:,NGٳ� *��8#��&��
C��15��5�	XX�P��1�¾� ӄs=��r�� &9%���K�K|֨��W.��!QG4V�T����N��Lp�֍���r5��Yg/\U�8����le�q�!���:ܑ�.;����S%�e�~f���Q��)~�q�pO~�i\'[7�F.ZNᒫ¶���h�)��#.o����~@�nϬﳹ������j�(`��k�qx����p��8fj5s�E��;sߍ�}���4�!�ߊ���l��p��B��ӈ�DŷpU5��r�;��8�5qJh<��O����^��Wo����P>B�-��p�o��կ^��%.-�>�ܜ��og�:M��r{����^�s��5���p��p<6m��Y�����b���֜0�N���k�W{�&7�o��J�k$���r��6:a��۵��b��+�<~�/J�p�̢�8�?Cm7pA7�#�o35��1�^>�/�k]]p-s����+�C�~t�ZY�p�w`i0�)U���+�D\!?1˥��oH�J=�)�&���Z�e%Xn���գ��%�nd"����%#�w����-:6���c|2@R��G'�`�UB��S�@���pN��3!(�cTs��8��[I����)��v\�#��k:|=�<X�!x�m|)��%�n<2HF�k	���/ٳ��
{��,��ǆ1�͢I�$���)���s.#�Y�У�۪w�G�\ #z{��$4��5�qO��.��v�a�� �4mz��kH�lC��4Z�5�N5	���R��'i�}T�ݍ"���b�g��)V1luGۓ�����3<�����.�?d"m�o����}�83��q)�)*8����L?�8���V��}8�����W48�vX�~��a�Y)�B݁x�Ak)��zͪ�pA��yǖ�+�0NJܸ(�E^&�XѪP@����p��"�1.���TVi-x��M��k{��b��F/*���.�צѬr�ۚS�'_ �?����6�4{�����H�!.g���dO��Be(V:!�P�D���CaR(-��$�5��w��1z�欫l����I�9v���nKjخ��"�����5xm���#�\ʒ�E81j.�CydxyTϛ[�>���4O���1�	a��5ڙ�C2���L�?1E��zm�-s�y6ƻy�]gHn�#ABتf�lʜ0s�sw/�w�`ij|TU�{�S�x=1]��e�(�"�����C$��P��0ˑV\0�+N y�K�)��}|t��f�I�a&[ Ass'y{�j���r˫x�? ��`�arR�2��L]���ɿ֩��[��eb����Q���5�h����/���WӍW����эOq��}���v<�,�e����⸌�,k��=�@9���	�sW)��QY���x��_[$�>ËS6-ƯsA�
�Z���B/��w<.�Zm {��+���UA]uL?�e<�^��޲b���t畐u��G����<b��<�`�5�D���z�"���ҙ�K��+� n��X�����\��+�ӴjW���R��F��@?�t�#Q7վ�����Y��$o�~�߱���'M8�V����ʯ7�9yMa�I��5��lԔ�1!�t�W����ڴ!�f��Utχv�o�yG�W�)��޽������Q�L�Y>�ɸ�21��n��T��
�^��	�}4�*��v"��T�ď�\5����'[�����b�%k􌀔^�D׃&�Ǣ$�%C#�R����+)����X�j%8J�������6��᫨�����@�t����>h��-։�I�Nv�S(��&��������i$<����k+%$�'������}�莂���)�:�п�+zIz҈ĉt�yu��E��ANl�&���z�_! �̕��ۓF�ܦ~ܺ*f��V%��\R�׋i�VQW�_�W��q�g7۲�[�W�>s��/H����-���Wyl`����D�W;�o�Z����oom��Ī����A����F���Yv(����O	�-������ �^��&���c����$�+��?��޺��":�}�6��꧱������M	s
��=�U9.@�c�~����et�N�	+���M=�U��O�x�7�G �;K���v�:��sm3y��`��h8?��:��I��z�\B�����X��ȳ�@� ��r�([��l�U�d[��}���&=�����6�:6��?kqQ��GҊ��.o��F	$�SZS�������.Kh��w��xY�>,k�������,���3���е��}"�O��J�'��0��;�F��K�J\Sl~4����+����`m�����
�ɪ���D�06��)o��u�Թ-%x����/5B�ԭ!�.�_%^���1�ܦ����6�r_��KT�G9A�M���ԥĮӫ��b>l
8��a�U{[Y  �<����Z0��U��{�X�F��+]��jEr�Y��0�I�Y�lk<��yyA[�x�[El-Ε	}Jp�n��+���/!ո��G)�}M�+̅��� af"���\�Wv�_����lgPwU��8ht��rq��n};":�b����,S����� �;t;|����gck+��t� ����K� r�&;�����yJ;Ws|����lo�f�B��s��h���!��fVf��vV[��h�.5�	��g���,������L{��3E�������Z|��gGQH�)`���y��W]�X��OC0b�!A�i Q��ml�<S����<�D��P�:@���{`�������;��9�����xd���en������$'��	=��E��`e;ؗ��]��n���`��O`M�O���Jc�C���՝�4gZ̄��nx�,���L�������������[ sy�������2���!v���J���p� ��|�*��0�������I��S���LT<}1�����Bs��8�\�i��C�{p��ʸ��G��U*��m�W�IvezC,>��^29:�M�����*���=}w�z�!QPlXp^�W~�yt[P���l¿IO��FI1���?>����&��u����QF�/��_]w���և���Œ�BF�d�J�������w��)��S|=�� �&e��׉8Ƭ`��	e�+s�9j\���,#�����_^�>��Ir�$��>2�U����>��Ǚ҈��t�T�Q8ޘ����[�(�^g�5��������0c����W����`��=N7^wX0e��r�G-�7�+Nԁ���}n����U��,h�:�/�;`�Z����m���r1>A���� Nc�[ᖖ#_��,S�q�Z�`L�P|��ۤ�;扼�kt�-��=t�`KV���y�w4u5�1'�������7�Ćd�
}P�$��Fq�_J9��H���U�}�;���O������0�T���V1Y-J6����`|�~y�!R2��#a�r�wͭӄ;��KaD���?���}�����jI����4���(�q^G1���F�O� ��K���oQ�e����F�o�z4��B��w��Wy�6�y�A�4P��S�S�idFuI��E���noR�G]��;��\(���?Գ�]U��ņŝ ���ݶ�U�;|¹W5EK����A��A�=
���9�|!�Ms�GO�"�e�.f�h��������3��UN�I �#�{%��#�7�}�:�HE^hzܵ"�Ɛ�,�#	�pB�͡]��}1�N+�@>섮�!Զڋ�V0��4�ի���A�{�eXHQq�Jl����/�J@DM��F�P1}���L��w�i��.���q�ȳ��%d�K�.U6�`���kH���& [q$X���u�r$�1LM:��:�����,&OpR雕�p�ё��ZRx �a�����$�e�?�b��\�#n&�P����b�V�Z�/�$a�p����̍��ɋ?Q���=Eʟ�Z�ǃgD)��K\ڿ�~w^	��-�Ӟ�XP�P7E�������0k�bԑ+�r�ai�̄���s��>.�[��2Ҡ��i`GO=�S�ƽ�g�=\�����-�`���Y�\/^�������I�A\uL��%
���zy4=f��E���T��]��@Ƙ\.�e��$�v�Kţ�]?(�l�n�<�c1�E�!���g�sܚ�a�y���s{aC.O�H�F3�kT(���C����s�MT�V�c��hH�O͜5�ʁ�r޲��y�8�dk�}Z��~��l5����5���`W�L���~C~O�ש(�p�4�_���&��(�{����)�u��u)�h�\n�)�y6<B�i�1 �[s����^�L2اf����t�!°�	ǎ���K8�E�:��;8��X����15ҹ�,�pٖ��`9�.�5#�.�j֙��9���1�]�8�W��2渗�i���7��1��F��~^\�� �"S�UD�h�,Q�ra�������JH�68]9��m��Lv/f%�E:��޺�yr9�� eJq^ڽ�����:Հ2*�G�{�4t�>���3��ఊ��9�}�����	o�t;3�#F����^˭qP28�;��&���&ڒ�Z�w�)Q��yxx4ݻ{�ʃ�B��,�|k$�0!��f����`�F�-Y�^^b 	H�v\�A�~�/}���E�������ƈc\-��{u�o�)������1��f��ꋛ��渴�~�#�	09B#6��	s�釁�� S���X�ʥ�8*�X��V�:R��L��|O׸�*ΈV��y��O@�	d�E헦 ���c�V7��x��meo�9����`ý<����/�ى�� ���N�M�4[��(x�>�z��h��%38�' ��A� E>�4�A�&�ş����`�=&�S�c[_A�顜6��7��o��6�h�葀d��^�aM~�C��s�Lu]�\ƁJ	OGR�
#EACP�̸���g#B�m�p׆̓osʌ`HL�x���o+���e��e2��/�F��%A ��(�-HX9�0�V��B@��J�Lb�t(�|����ğ��T��Lt��y�Cq��C�l]���מ��:����Z�I���ٹ�x��z�����'+5�i�����7"S�1���� 
ۨ�d���g[IeUdId|��Ύ�-�X|�F��8���1��y5c�����L=�(+,�ê�&�{����z����'����k*Ӡ�3b�ۗlt��A-�n�6�X��ǎ���r�����f�q�A��=�U�ĀI�����6=�nY��}��c�v�}f�ѵ��?�n!��,3rY$���f�6~"���+�y�\i�_>�$�<�о��s&�;5,F�K]XPk���C�2���ʧ�o�Uwd,U�G\�Y���ټs������0�g�!n �g�\!���u0`��ǁCMd(�6�l�w�t��D�9���~����L�傥@� p�w�_��Nɇ;v�����H*��Y99VT���k�J�""��F,�;I�M����rU4� ���N[��@�B�2ԂJ���(�
�x���Y�8��z�;��@mT��[�V�8�L
�߆��R]X�<��R��i�>,��~�|�����Z�Pkʘnٗ�Q R��?��ƫ
�s����Iv���jل��n�w�M?���x�V���]��WJā�.�@�*�<	�J���-O������p{g(V�
E�W��S��`���-%�����*�X��) ��h8�U�o�j��4�3T :Y�f�yA*���z|nQXN��k3��΢�_����U������ki:����t�It���\㮥~��M�ښښ��/�s�2(���	FvUYs�n���l)���lJ�³ġ��A�g�ja�ʏ���4aX��b~W�o���g���K�2D����[�g��>�qs�WaK��W�@��Y齺j$����;?1��ޕ�G�����r���a�MQ�F�c�����o�t� ���ٞ�fd��iE�Wxzǁ���P�"�ٮ������g0�{|Fn#&�jv��3��1���!�����˃VM��� Q��d�P�?�AOp�̺N����	�l������j֋�rti��ĒN�փyt������G�'���,M�a!kԥH�aa䡹���}d�T��^Z�Q�5���������<�t��녱����%H)�.c�4�a?��¸`6I*�z7���֐x˄����S7�V+F��'�P��D{�l�Ù�T:�� N)I��_(��()Ѽ�;�(f�D@��F�����8�����g�y\�8�����z���Q+Ҽ���J�1�c��_�}������t�s�LgxKG���[&;�u��<��U��A5�r|��D�v��Do�?��l���y5�LiT�t���r�8ܽ�8��](6w�삮q`3h{�(���^CoW��İ�bx�P_o��Z����7o	ǻ4D؄���QSv�t��I�\KM�Ύ-�<.zD�m-U�|��ޠ ����1 �Zi+�K�!��F4������-F���e0���T�eF))[�S?)��曁Q�>�V�I�;k
Ʒ-��B��E��I�fچ�VNf/'�����ܴ�j[�'R4)�`��I�h�����(��\*M�Xq�N��rۉ�״����#σ�D����>�ߕD�(�q�4f�4~f7޲�R�3� ���^�u�gY��N�$�^�6���.D�DE��C�T毬^�@�{�LA\xoU�dz[���8K�F���Xz�� ��Ȯk�M�2Պ{�Y_�73kK	XH��yEw����d�ɜZ�#�����yx�.9��b���t�oϡ9X�_�>t!*���>����ЧںeLT�s�)͹��H���_��O	|� |���wR�Q$yMFү��0�
GnJ��{���Q֧6�ʘ!p��ڄ'��f����1��.9Ԏ��E�v��I�=�!��J�R>3��g�2��2���[�6��}Yݳ"�p�rS�1|�<��fϞ��/pĆZ��çtB� g�A���q�uЄ��K��
8ù��zۻV��yF��cP�5�.�7]����'榄l">((|�s'��I��^b���-�W��Q� =	� q**��wW���d�g7W�Z9ڔ��o��d�36;���S�\ë+�r��uޓ!���'���G?M�CO�Y`�R������Rpd�2�aȫ����;�?���7;�0N���1���]j�l���F���S�8�"��z��b��C��RG
��'�
�:&���J군V��h�!��\K��+���?�&�d�ʙ������`ީ�;{p��4�Z@r�N��\j����C�N[I�C�����T�&��#l`GjA��_��~_���F\'�m��ƃ�,���ƥ������n,8n�� ���L�aɩ��H�w,^�B����[��Q�(�hgN�g�Iז���D�����C����En;�s��*��@����  ۿN��C����T�%�(蔖a�de+壭��q�ޫU^ذ@�=fADV�� �o�f�`�T�qb>9{|�kG���A�.�I�Ȭ�L	��OtmOT=�l������#�W�cjb�25?�5�1
���S|��uo��ʠ��2x�ȑbC0�x���ïI:P�����x�|-����d�T�0짙� �|��#K���IV4G	�j_��.n��c�Q8��Cx��ʸ
p,kS$�[g�j�@�'�`y��s�IBD+��ףX�#Ip��Ey�ee�7��aw�����5�f6�M��i���%p��_��u�p�������h]�ٙ=m[���1J:�o����:�i�L��H�BϤ�B���m)�g$����`<T��b���ݼ�đ�Iמ_*X�"U�����e:KM�~\1�/���O�|Y
�m[�c�U,(�Vl棜m��g�&�*��ޚ"ˑ�p���m�d���a"�{i���W�7��O,���w
Gd�_��7i���DæU	�UJ@[3HHi�8ft8C1�)E�)/����&�R���(�yw�q6PZ�iۣ<e�I�>�W�/VC_)�� ���w��_��+&9e�@YA�� n�f�c�'<��.�^��y�}&O&(G�'L�g���>v�֭��|)r�O\J�t�Ձ���%��bi�)��qg�m���}g��h���Ce�:�l�����i����}P����)���.��[�U�d�8$g���C˾�[=�	Ky�w6�׉{Uzy��;zDfQ�?W���=�NR��ů������Һ�r�3In��|��*�9���V)��RG8%N;�D�rl]#����"73Fo��'��ybɕ;���+���Ua�t�T�09�����>��4�|��p�2�:�n��38��>	�l�����6��y���x�d�u6��f��Oh��S�� �����+���q��bd�<����6��x�<|��7{�+6�[� �,�
���|�v�#��RF�!���a��-���Fa��۷|�M/KCOi��EU�T�aR��&����������d�?X���@X@c�?/��r`(fH4����lݗ��5�~xkt����aŸ؂�3B���MD3yUsrr��˶��� �Ӊd2ߟ+2���3N;���~Z�+�3��oݠ̇��.M�|�J9��
����X��;�L��9Hk���H�j�0�,�|w�ǈ��d"�
nv�s�]_���p�RJ������ְ�U�,�%>�@R���ӑ�n�Vo\���z�f�,�����Q�H4#Y��۳_��u]�'���9�ᩜ���q��$�_�i�U��SP�#U�8	U,
<�+��֨�$�}�'�Xx��MJ�N�������	,��C�q|�2;�I��KA2"�.@�T�?#��1�?�_��!2Ď!`ȼʺse��d����>�xq�A1�~ռ�X��r�wp�(=�X�:����"7����X�kJ����;�U]�:������g��
��-s�<}Z�*'�S'��,��|,�]y��8�A�ٰ�֩�!�^��9���.�`�k6p�{,ps�B�{�yc~vj�z�u|y f���P��Y�ڿ <�r�#G6�t`:ݜn���Z?�爹��H�=ڛq��@�H�9L�vM���z`�����~|��kڕh���'g[,p������vɷ|#넼����C���3)��F(>�(��%�Ƈ�&�_{�����2���b��'x~����O	 _𣣢���ܜ�4� |DD�2��sJ�!A��4�p�F1�o����#u.�mh�br�൯3�5}�c��u�r��0�H?��v�Z	�.�*����v�[�qwu����(�Oey��o��9^̟�^^]i�����I��SK_$ʫ:0���8��9ӑ����k[�"�=&�%��A˃X�YW����ƜG4l�0'��>����t<�$H�uJA6�,����c���[�g�����gT�����Q;+K*�\��!G�A����\���s��[� ð2c<8N�_���9�N�'�N|�%#�4d�󷆱�\}ɰ��� �R����K��6�ֹ.��-��/��J^,��L�l	X�
D���)�����@����b�k���ɨ�#�z|g�'=����-h���GV�PN
�`p�wj�B5ZzT�i���s>��f�6��#�o'�H�G��_�B)��#1�i�ˀ�v|�[��D��-ӏ�g���\�H�Z�s��}e�CQ���l���.I��u�s�2�6��c���E��'[�>���gS�(S|$^K��H��P�qG�i�X���<o]"�B�Od���I��Io}����)@]�̙�8m1I4aOC��!"�ؔ6���� ��]�2P jl#�1�1�`�W�S�l��S�_�,Zmo>����Ȉ���"V����`@���)v�D�08o9TٯaPO�p���{`2��N��Jw�S�k���C9���Co��/�+3݇8X�%5���H�����ӿ5���"H��!}3=�q�S'�3���ൢ��mX�&�9��׋qe.@�Hz���&n׮��	 ��S�}��K?a�7-Fch ��n����b��,^�/����A꜇���S*��8hX�}pF~�9���!e�/���!#Ո����<�=�^��ۆ)3�\n�r��Wr��kh|-�Ί�.6���s\I:�Z��8�J���%aK�L|~khH�nV�r9HV�PX����#�?C�\A}��2d3�Y9�k�V K���K9��%���dm�QY}��m7�k,E�2:M�yٹB��g�PX_��Ё�9�=v��Į�|��
�!-��p�/a)vJ�ͺv�u�X`�ĲH��Z�xm�d�<�߿��/{�� �q�
=�}(�<|���O��Sf)�Q�ܜ�]�w��][����ˢ���?���� A�$8�0��d&s�+B�K�͖� [{V�ŀ�}�{�ZM˼����L�;�C��Q}�8vNP)kW�qo#���+6K�/)n Ղ�\=��W!�d�������ӝƋ�r�3|i<�"\:-֖�#��s��_`J���#n����h�V�tr�C�1Α�Y��#��Ӥ�pv��F��vVB� E��YM-'�q[ԛav���`Ӥu��L�Zo����zg�����a�	�T���̃t%������\70�]'��jn��/u��D��mԪ4RW�u�/�w�zT��*���68����
cFp	"�G�L�7%�\�<]M��9��B3r�Y���O�G7Fg"=p��f/�	ΩSPq�����>�i;������]~@h��5WMm���0큐���K�*L�"Y ��t�VJR�p /�a��2�-��A8B)E�{����C^ ��&>�l�؜��]&.��h�{Y0z"�֩�e��7� n��F�����e������<^�8����Վ�u�q�?�Ub����]� *��5�(��k;���gmOA������B�h_8�׳@ �d��Yv����Y]���������-&Z�"��������s3>�+��K�:(�0��
�v�t����ԀH���G���6��R���ĺ}�,e~0��)^���D�q�[��������a����ˉ�Ӛ��8Q�Pqq�j.���!�22��DhE� ϑa��'��X2!��i�E�5E���2�*v��"K˟F��{v~<�crɷ}��Qխ�� |�"����:@��'�>�z:?S�,��|{���͍���Ce�*����W� /�jƻ��o�É���%�lm��E��`kYKJ%t���I��� u�wx�s��tU�Be�m����d2�pw��ﶋB�v�ˊ��"v� ���������	�6Jr)���nAd��c�a����+�c��j��:�i`�󏠇"��1�!���myO�t�"%&�6���,��8.�N=E����P�Av�3S���f��	1�!��[Ͳ/F1���7�"��.A\:��k�٤�|�m�(K���2�&����m�����HԾ����Cݻ��aj�ﭧ�`<��2K7���_��f~���jS�c$�2$2�ߵ���偔%V`f�,�tA1��|e0��:�����$�'^��\z\)����HаD� ����t	����
��5��|~8~���Xz�������Vv^K���K�.J�bì�����Zp��jp�h:�4�qʛ�3q���I�|���{���K�W���l�6lVL�n�o����~Z�I�2D�y�S������gg\�	�w�NyL5�6��^ g��1��Mm���-�|z`��Zw2f�²g����,��#3���(?JD\-�6A��t4��sͷ�ӈpM��q?{���(�%ָs��kg�����͹!�Śp�;Y}J���l
��9&1%����T�ׄ�����M[�}k3��Xu[mV��53�`� e���+|m_��)Y��%��A����
�����4�n8+��m B����Qn�^p���b*I���O� �1�Ok�}�������u�G�|�͎zݻv���l��.2!��b&䜻	��7X��$���y��D���P���Av=8�9�u�f
�E�6:Iu���.��jJ�<�)��W����D�ŋ9��~�TZ�<%����U��oҰ�y �m�XT����1nV�ȶ�s��x��>�� �q����?Nv?�@�3aGS/�V,Wm�솱g�'F}"�$,jM�����*�ge���63�ge��a���a_M�@�u�+.�u/D`]pKl�}d��f���Ǣk� ��\��ܿ)+�������_R����f���߀��3���I_������2��cF�{��A�!@�|L�J6K3��ˊ��Pq��R�\�	4R-��Â}1i�u�&'n�-�b���m�!��8e�He�j�A��?T�2��1|�2k�f�q+�ۊ�\i�=�6�c+��ȋy�[��U�Ά4�Fgp����xq����2�Q�H�@?%��#�F\G4��,A�{�c�u�x���r��D���a�wo��JG�jP�XW{���
�y	B���å*���4�2�vo����j�f���sO����TR&�*�0�Hѿ�CVb[.�z��t(�-f�9S����O���zhɧ�D�k��K��x����U�2]Sl��o�m����f��2ߍ�O_� dp�mo���$2������L���"�����k#�0C���`63uS����ywDx��kf�,�\�,G��:>��T�����c\
�gG�Zx	ש�l�C��4�sc]�1Bbb�k���Zt��X�7I�8+��㋗�33���V��h�FY�A*��B�q��O���F��b�X�MA)�
�O�����"L$}��D_�ȃ�r�rO�����E>=�j:�ډI����4���{����Q?��^�?Q�c6t�jR��t�aW��상�<�C��Px'?Y�,Z����b?`��RS��7�u�
�1�����i��1k�|�P�]�/-��SMG' �����b��!�=MiM7Ok�nN�*���q*J6B"*]�m�}Ν�n`�*@5T��!0���]J��TC�x)�D�H�E�B�V(г��2�.K +�.����/
 ~���!倷����C	݂fΏ��%�v8ֽ?�wa2�T�.�+M_�i��ό���O=�V�A��1�*�o��9X��yჴ����{���"�ٛ%�ωkVr�s��I�^���3��nXas��S�\0�NB�2�m� U���D���C��Q�<����G[��@j��>��=,�vq��HyCk�лx�.�9��D����;�D�Uџ/�#�-��us����=Ҧ��/����p)���9��ǳ���r��qR��=���R�W��nP?�-�#� �����)dFQ|�	��)9"�l�X��"t%��P����<�|B�վ`�&r����8��������n�ZVGC�$�����i������'e�[+ig��}�F�I��o5\�v7e{&���<�v���VCX *V|�I|o��ǩn�(��b�T'1L8b�w��������6o�FR���.��utW�4��֖ۜ�Mnը��U��h�>�(��8�q�@��{��=f����l.������1;2��U��G�|+��<Y��PS�4��(T���5�O;J �F�+I$�G{yjՂ0�=`����S��ciş��5SOO�;�E�@eu�z�v�f�e9��v�F]��1�>�9]�A9�E���I 2�����M6JV��R(@l���h����������lW^�uCh�� �H��Z��7u Ҁľ=�B~�!�<�X��B.���W���������S%Jt�Z�h  ��'D�A5�߼�mX�J;1>>����K�dZtj��K�u�����c�q2$Q�ٍ��'�ǻB�ʳ6�JL%��#���X���pī�Oi��n�������7�A���#]�0�!�q�/�Y�"3�d+wj�z$)�6(t�G���L��Sj�K�(XP4}Y,	*���o2'���蕊<I�B�m�{�)�8γ��jH2�4��� |>���y=j�=�Ӣ�v�C��J���a�\�`�����D�N���Dp���q9� �!�U�� �1D��g����_]5��> ����7���v�p#��8,+�/��~����s*�V�3Ɵ�W�!�ǵ@_p�"b����	����n`N�jJ���!���	tT�	J��{��r�\�0B7l[͛	��S2�a����0kg����gQ<T��иT���H���H#�	�,x��`�P .h/P��2E��n�(11��<��c��}�q}#K��DV���$/�5@�b`r��E�DT���f��;�|n�:	�=D�����Q����o��M�f���;��:�p�!��̸tQ�b�j�U+9�f��F���CkMZ�,���vxL�Gin�fD��C)�p6n��(%:�о����Ѩ�����Cd2��N�V�&/�����'ڏ7�����B�k�cs��֝�����?����!���A�Z��%#9փ�}V)�R`�H����t���3I����J-��@��Y��P`��Jb+D8�Ǹ�x��@j�,�ql��� �m��>XY�����*����5:���N�>�Lv>���_#�d��,�J%�f�Pv�;��guk��&k���ʍYQ��x������¦�����+��(���.�T���_��$L3��;C��N4~:'�&�ܐO5]��e&�СQ��[��@+%�=F��N������ί�_�CΣ�iw@f4|� �`���BH1��]����"c2�9,)��Ү;1a��s�����k`~f�)R����#H�����}(?'Ԗ(�Ũ��1|��Yߓ[)�Og��'��h>谥9g5��G0C�IQ�ɔ�����չcd��8σ9��50��X�7V���dm
�W�E	�_������|� ����K�#-�Z�l}�Q��pi���[�c�'�����$Vk|�ǉLu�)U鹮�~6M=�����ZF7�j��K5�O��fh�.ʶ,�z��2�4���y�d]-�W��^��m��$,~��k���yudM'�Z�M���1��N��̍5W�A$���T=��2�L_#UZ��h�*R4T�F�;�"��d�\�1�n�'����1's'e�fc��[h�6��,ʔ��p�cѵ̨��S�+�L!������/��YK��� ��ł֦����
@� 3͐���J�O���?�;4l�%���#0Z����Cw9=V	$$�� �3j1�*y`&���=Rv����,�������A��jo"�-4�2��dx�A{�"��U`��_7�Ʃ�_�^��r���c��p�7s3n-��w��$�HY2V5�P��5;+�_�3!�A��/q�\I~�:�<[�I*�����s6�[���~�͙�)&����1��SL������5���^��S�Wƫ�E���fU�*Fby���Q3vf��6��_?Ze��E�sHv�%E(�iv{�C��CZ��'�D�@J�uj�}:�aqV���$3����#�~�Y��2�<|۩��)d���q�JGؾ����qy=�]<�V��f����͙˥ax&Q���Y.q0�ϻ9�싏)�����f;t�z_~�サ	[�-�6=�"}�m�>�Fv:BZ6�OۅA��E�����8 �&�(X�/�Mq�?���xC������q)�~LQǥ�}��񮿜	|�GN�|�ֹ�;V\(�(���R����Πh� �\ W@<�~�7F!�U�#��Arv>��<�8�Q���A&r��bA[~gZ9�w��_O��i�i�^���p�r�|�)�ufҰ���� j��$4̍D��99"�`&d��{�2`������坫���5`&��oF�c��7#Gk޷�'n(���R넞���s �7	;7<�:�F�}N�J&Y
�JV¶,qd�֮l��d ��ٛf�dw�t�\2o���uWR��]2)���pm��r�P�>�ʫ+���v��F�uΗcU(o�I�έ�����I���u�ݘ�ZK���Y4� �i����F�S8��'CJ�nU��]����9����	��Wi����
���z�'<�}�O�n��e������v
�����Y������+a��d��hr��� )3�r��M���]\�Cg)���}a��bʹl�R^G��b���W"<98[���Gg�`�d��L<Fe����v/"�4�t1oV˃���byR�/�~��,��he����MW�{��b�}KO���d�g����200gZ`�5c�F�r����O�sؐ(��&�3�Ԣ��?�y��l���l�ER`��o�K�猞����h�߱}����ݝɞ�[�����Pl0� ;�ͽ</�s{毝�7,c ��-]�:�3����4��Ԗ2,-��v�*y���!�7�G�Z�l�aE�ߨ(P��Z��۸��)
���I��K�A�Gk�9��OU��"��`C�� ��'�-&���� F�.�0�P�ج�w�$ �b��?�]+=�x��x�L;��q�)�DhR��'��j�-��m��zE�5�8����c"�F�yG�������u���x#�hx�l��
v{�?���L0�T�҇��fɴ!�J��O�	����7��ț��[�����]�_e@z50wOP4�]�yy��܄��7���`+��9����Wچ
�ke�p����F}�ɋ�wD�X>�l�v,��ՠV�����̇��B4p9�i�G�� ���
k��ُ��q-FWc�ζ����!���S�l�忠�)br�M<������l�h�1�tZ�p4�E`�A���-�UP��I��OO*��REkm�O��g���l.� ���n(|O�*�2R=�"t�$ ��C�v���
�$r�aJ���>$7����k�nz�����0��)\ �<�Ԡ��.s�as�]��6�r�b�~��_h�� ��ei����T���:�@1��03�]5�Ǟ�.+o���O��*Ky��1�!=��
��x��y�G�\F�ЏM6Z����5�ѵ&C��r�g��=��\'?v)�-1Ir������K���5ŷ7$T��|f�s*���z��5Fd���\렣$��JC=�{ݍ�M|��+��QDC���yxa���%ψ�2r��.��h�](���z���*��Vi*#d�~źi3	�6`��w����f�����u��V߮~�W.(~���^
JLպ�KW_|��f���Z{�ݐ��R��g=���\�Jd0WV��:��C���ɰ���ގX� ���4B� {��h4ΰRZU�$��@��/�*��6t��44���iɿ�V�w�5&=���2'��}Hh���Y�j���5]��+��F�p�j����4��kl�i��Pz�!���N�{[�d�#nW��@-�yXow���/��-�B;�.yb�w��Lّ�ʞ�`~kzX��c��������&�L_��e��m�pPënr�P�0��w�L�B�*/`�	L�����	<��o���PP���-;b��C���8�伉q	q�0#" ]�%����p7+EyyR�5p4#T�k�@`������/âN���I��y�#�\(_�vi�uY& ޾�MS�h�G��:�.�U�k��q�dF�*�. �k0��״ߨڌc	7j`_�/M���uO�����m�'$�Oo* ��B1|��5����>�@�ɪ����Wy�<i�I�cg	��-f�HGd� ٜxk�hу&6զ�^��4�U�@R����@�u��#23f�;j9��sg�� �9Ա��ɸ�����P��w��Up>����Ķ&�|~@	Sԓ�8�8�1 �
c��I4�ʥŠu��7��Z�K.�蹖5`�@3E�}|���l�:l��ΦI�䇈����_ծ�m�d
�oJ9;5E�`=$�	 �֙�:�Ε�,H�W^� lt˦�fUF�O�In����G��(���*'��I���˲���_q��h+�>�ON������#�$�a{� �&� q���<�TT�̽�V��CڡץP�����q>�Mv{P��`�t��5<�sq�ۏ�g�
�Dzѽ��KfK��)�۔Z�m�}�=[�0�z�H�)�m��@b��oM��.��6��k� �[��6W���z.!L�Σ��W�(�ǹ��Ie`G˨<}O�#�ʂC#���G$�>���n}������`��>|E�;q�Zf�c#-A���Շ[W�ɦ��ˎ�jV�n 	�7]�4n$��,�2�����fFn2(X����&D1�x%��]P��6FA�f�^���\��w���۳���%b�&ik0U@����n�ߑ�����fʙέ;��Ҩr�Y��ݪvD�p;%���3�Y&;�|J>kZ��V�	x�]�yr�����;Y�/�3S�oA��ז&rus�5u�-Ja�s��5��:vg'6˷6 �k��A=��@s���T�X8)?i�e>�2%h\]D�KSķ��_}�lJ��|�2~�l��ԋ+� k��p��K!l������#@�Uxq��V�۽���)�.M�~�i�L�"��7��I m�A��c���q��N<�!�J��f����+��l�T�^r�45���̱����v�$!��N�N<�%���d+��v�5y�z{��A�����<��W��@��_z i'������5\�H��o��J��V]�8H������>��Z;6�@V��$ky��5����Q�����ypi�3~���rc�3�S�$�'��Xr9��m��fAoC�����:��	C�X�d~�.�:�rtYߴ^�Ŷ�P�&��\�5)��S�]Үuu����858��La�F�a�?���n��TR̤���U���?"�T�'Z���q$�іV��p�/�(�V%m]T_T���z�����������z�G������.�~@W�4���0��#H�������ڰ>�ɰ��m�V�RBʌ�?W+t�x
�N�*��t�������Vl�%]R�kG�0����x���&{t��$��=���q$�T(�oX��o� S���X9�+~e-JW%�Zb�Ș˲c��x���3Z�]�+��ez�.��N� N}�E^@.mQ�Ua�y
oS�u���z	�������[�>i��n�r��o�FY@,�h�b�0Q�n�]8�_$�#0Ʃ��SI�� ٽiĮ.wK�YZ���`��噰X/N��0y�Hք�د���L��H��j�>>d�_C�-e�p�|Yj�]�j��6;����zZ�%�QJ���A�Ȯ����$��?�O��H��GS�6I��kv��N�[�_D v���m�8�6$��1]a2P��j5�a5�ޙ��/H�\G�K�tf�3�K]�Qcc����/ԍQ��E���#��IA?��%B-�H�ף\�d�"�Q�}̥6�㿨S��}��2��6tv�V��眩�0J����djz�ON*bm%l��!��F�n�a�iy�H�'8S���#�}�4JxާT� ��� ���'"��F�?���b.1����g�����|<y�^D�$�1�gk���r�����4���Ո�)��]�H9X�.���0��P F ~���Qcu �����Ʉ��nc����:��xa�ڛ��L�/j��M_��'�&�J���7�c��Δ�e[cw��k�ݷ듰IIdapO���	lQ��<+7��E��TN��`s�Ωx_âweq�c�[��
�b�����Z!�PC�K���h���p�@͡���'p���W$jh!��G'mm�rm�YU�Y�e
�kwox����[	��\rf޾�s�/i�ǭ߶�i����A^��8���d�j�|�<_zQ�7��.�b�����V��g�z��s������ٌT�W�Ak�2=9�=ϧ������' �.�Z�En�K~��6���}��ڢ��R�ь}�۴�AW䞌7ʘ0ҴZs��]�+�1t �|����˯�pUO�p�� (�>��[>άc���c�dFd(�@�X><� ���n_�7����y��®�����[maY���hx{�W��$����Ѻ�|�}M�9�#�^}�bH�p �	.�D�J�A�6C|eVD��\�'�rG�q|bn�(���3�)��N4cj�w�媴گ���{ǫ�=�f�8|��9C��^�Mi;�MĻS�<��3m6����M*0��b��0��]��*O]Y4<�E���97jC�^a|�� ��O�l�̐�fo����9R��E�_z�y�}�
����N/I_ 
r{���tQ�t	�L0�z����Kc�gb��/"C�^ALW�;��3���ek�J�ҍJd.4��z7E����N�������ݍ�o8��w��Z�d&�C(�&-�*�wK�j/���3���D��4�וq!G�L��I0���Vc'Fy2�r"�-����7�_f>�>�^���X��x�?����ؔ 7I.lB�!o�α�=�����n*hoqa߭e&Mv���|����&��=r�J�f��%���M�w/��&Ǌ9�gD�Vy��n<�D����#8���H>v|�p t$&�+3�JU�B)��(�2��&�����,o�L���lo�zmC�\׫j���X�q�r!,�(.'�\��}����m�%ڸ�ʺ5[��h[C[���e�sYx�H2����A��SruN��:�۟����D��óAu�'~'9M%��߃���2ߖ�U���������en%x*0�ZT�K�Q�V�F]�ߪ%))I��& ��j܄l��#3t����Q��{0�p�/W�P�� G�酚�g�wV� �d���w�ך\���.���{���S�v���m�=��+�,ln���!~��2t�"7��D�:Pb�W�4�%�-���p�q`j�dK�N�2�A�S[<�Ru�H��	%^k5�qCY���9#�Yja,���C��hhN|�e��A�-�s]��5T��̐���I�-���ufz]>h�Aw��͌g4z�l��޹�� �}�ƄU&�5�W�o���
���r13��:s㵵UHC�Z��	@��J\%,I����χ��E��.����l����OBa�Ҋ�l���)m.b˗A/�C+ǈcr�m֒d���;��7���L|ײm��7��ɽ�p�u���dn�m����=�>�S��z��G�ζ�;��r���F�D�o3m����8�IW�BGE"����/�f5oQ�c%[�[<�r�ޢ>e�L����í߈���6J��wLj������{���1зX)wR��Y3D�.�<�����N��n�4�<!�e�:�[ErxTS 2(��E���ޭ�����;tV�wj���i���@0���u�#kp��H$�ʞq���v���Z� ^%0�ЫS�� ~��1�W�=��@E8��[�������6�=gjF�Ñ�s9w�]ɻW��{�ܦ�|�I'�1��#l�,��H��yV�S��-Q�RJ��d�C���?��b�s*�71���-��uQ��g�rr�QK�QPRSg\�D�q�r�]bonR�ث���#k|�52��]��5�*�]�����z�&��t�Nb����Y׺�gۮ��}��!��J��y̳�Λ�y���N���-�S��v��`��\����A�!3�Z�Hp;�7;��+�W��]�t�oZ�S��!1�u�Yg���)+>�x$���2��\÷���-�O�Ǔ��ءL�~6��VƖiGZj��t!�1��k��G!X�n��;O�G8ƔJ�U�=��&���	���W,���SaYΉɿo�"��Y��>ާ����
��]��1J��3߭�Ȭ� ��u�1��[���E������Q���v9#�ѱ����iҐ�=د)���ow�!�]�n���gõ,�B����>��LV���k+��WТT*�d��o
w!N!<���<�(��|uh�Z�)/V��E�V7 ׃�q|���G����Rյ�I�/��Rs�&�����taȊ?��`M䔊۫Gz,�y�|�!�7-���+^YgO"n���7��/4�w�� E�Y-P�cV	z�;yN�'���P+���98K�y�n������+��*dG|�w���W(� ��8�K]A!3p�� vV���̰��ݥ���'��6i^|9�ͳ5zz^F�p��XZ�yj)c�׍�@�/YƬ�:�Yx�ABL�?�b*j�_�"m�ѵ��62��!/��5��D���A�T��qԨ�B�%`J�`X�@6T�0��� h����>�s�5�H������F�sE�/LY������F0𓱶����,�@�tt'tm�O^��Ó��xM���V�od�P^���{rU�	NQ��^����T��v@��9)���<'4��#�������ř�,���ŝ�\*μ�|�Aw�}�7�(�*�׈<���5� ���u�N��pX>��� Ľtϊ���%�1�[�!pyRa������W72X��pN�o�-y$���v�?Gw#[�Z��.I_�R�z�sy�"p��V5���e�s�p7Cia'�!/{m��h�MA#��C�?CM��I�Y?�B����w��j����Ϗ�s�I�pg֚������.f7M���0���)�]��	}���~�"t�DG�"kN:[ϒ�xT���'u���	ǄU����9�4��	����k��Q$���l΁ҟ76���6�]v�S��_�x���{ؖ��p��t�@�ֿ�ܔ6KݙY;�Z!�p��ypr�W�9��\�����5ɍ��;�"Yb>���:�0�k.��0��=�<J҈�^*8|5���G���({�3�I�^	幀6k�;�&x���f%��ȓx����Rm���A�L��1�a��a���}��V���6
�ZE�]�7⚟S���k�j���@ɝ���pX,N:˵c�J<4}�d��kT4���9�F��\E�=�Ŏa���;r�g?[�u�.����Џ�v��:�"y�������ːh��/��Lv�_�D^Cu�|��%%t��l��i������f�j^I�o���UV�7�4�ѹ�7�P��N6&�f {�TZ[^��3�{u�[�b�n0�� %��NnD�p�#UQ��'��6R��"K9-��Nl��������j�匒s
}w�'�۵rD�S"r�V�&��%߈�(������������g���l̕�*71	��U�6���E���B���U�
9d�p��F|�l�II�7֊P`�m�P�T���;أ3h���d$ �V�(ҟ���K)^#���^Ł<�FT�ځ�����u�������ol,�Į�4�n��U���0�2�����onu�P��&eM�.�7�x6尬�!9��T9�Rݶ�~����ю�Q���P��Ց&�#e���I�I��8��E���B�/���D��x���\�%��'�36�"Y�S��Pf���})U�ĺ4�R4 U���@��|pt�z��Ϟ����$%���0���'�Ʒ�h��2��0=z�����[8i���! Ub�;��������m�V#�fL(�x{M�`�P�X���Jf�Ҙ��|`:�kW;V"���YE��s��h���@p�����:/Ƒ�<5?/���4��������*	����p-믝(��_�8�\j�m�ۃw����W*g���,px��0BO60a"���d�װ�D����
�G-����v}҄����ő�H�VyrW�W��[��+�vÔ�������=0�$�%7Z�UY�m��@��H`qN�l�C�;M��hu芘k�x,��4���7��R��qWípO:�q�L��hr����V�_)=F6����욾N���Xۊ��;q6�
���,�q�L�=��u�Mu^y��:- ��&��Q�j�s�?9ܐ�X��*	����{�{����MqY`;�h�io�!�2�� /{��`|'�*�N�q9 =��'����~�IN���i��&��+�;�> ��e��$T��O���`�6���en�������2��i�)����B�IxYBb���u���	A��m�3��L�oJ޿Zx��u<����/\=��9, A�3�9v���\�<u,�l�;� �#$t��B�P�^�,��V4��9q~�,��˰|����x��y�R�����̋�Ͽ_�� ����lIC��x��"�+b6�-��K�?2
��X�Y�\C��kG/QkuQK\Bf*b&fv����u�8{��q�y�%V�!a���?���R����j2d����L��d�T�H;1ֲ��I�	�6b���ordu��Q�����Y��@�/�/�ʃ�n?��7�^\:�)L��5�@�g�5�T���"�,8�﨓wÁ��'���ZAzx�o�G�ӹ&�6�*,BY��xQ��V��.���wEj-��(�F&Q�ܛ!s��|/U�~��4���'����&,ZB#2%W�|&�yR�D�h��=i���|�S����Ѷ���V6�)��v�dR����L�8i�=�^��{TꀎM���s�K%����z�&}>Եx�ph)�UmĢ	Ԁ���X�y�9` G�$��7T�D�����6%�IO�1�ʃįH,�pHi2����B#u�~��O���2J2q�tFw��l2�{����4�K�j�^���P%��+'
r`��7+Y�й�0?dI�JЅ�'}�:))2p<�����O�_(r��W��OV��l`5l��{ƺ���=��s����R&O�I���V�5�a2���J-��R�d�l�"�|��-�9�2�d�zv��8Iju4����
����-#A�vQAgq�E%���I����["	Ɍ��v�d�����eĮ񩃕�O��6����`̮�c�d)c��S|��i@�<XZ����qn�H)�����H��}���"	��џ$�y6���f\�I{��P�qN����.C�EcbF�p�*��������M�� w� '�.�]R^�7��'u��yKs�vvfhC�Q?c3^�	��Rh��m���*\W�Y"�M��+�]�ù�1�4����NJ�7��t��f|7��/1vz�����>����rDM��8J�b��N�t�m����=Ze�GS�� ���룧��IL��|d``Ɨ'�ԯ)'���X�L��M ��V�DT�l.o ��.�����6�hϺ'�GE�M}�ڨ�{i)| a�b�bcЭnO@M�D%��2�~17�⽸�߼f]W{e�3�I����AA��[C�}��r���j2�xsւ1ul�e�߱������\�{'D���I�jĳ$cƙ0��ԟ@۝�a���賌���k{�g�@�A%��߈ha������eA\�I�2r �DШ?Nlpz#�᠇���D�q����m���)�]�[|(D�g��?o�e/n�cnD�/X��C�q�.�s7�3�o��R��=-�M�X	�@�A/�`��:]ٷ*8`�'X�Y1�� R�ݖLꃍ�\�l3�?�:bD��#�w6� ���]���褥�e��b�`,5X�]3��|����ҍEg��;���`��4����T���~d3JN���rT	��(#��n�0�c8fsY���Һ�y5�>K��ҌʊsH'�E�����y}ѕ[����;��>&��]���Fz���;�)eOy��]g<�q�ވ�;(J��PnL#
��F2�I6:t�iL#%�Ve�Yx"����^��2>��Y�=��O�����?�&H�J��*���8�C��`��^)F��'%���L���2�o��1���f�^xvl��I�mt(\�Ő��-�(�y'EĚ��oFJ�0�A�3�\��Z})�::�%����h^�V�R�(����xf�9-;=m��\��k5�J����]���:e�
������<� 
HuM�N!�%��q�KHRY�[%_�ȫ5�-l'�Y*��p�� ,��Sڻ�8�e��J�0E�]R�\WJ��	&)�U���=���H�5$m)����^n[�k_/1��O��SK&�%#B;�iM(����0j���ϗ��� N��%�l�f���AD���׈�!�9F�^��_���������^.���� ����ĉa�]�F�����T�b��@m�I�N_��A�y�y\*�=B�1�.ˋ������+T���x`7����'�e�c��c�Y���}����6Ҫ��~�L�k�@��j�R���ZX���K�HJ��P �u&���w�T:m�`��"_pxD�K�6�g�� �2���e�Xf�1�B��ʳ� *U��q�o�SL�z�����-�7�認�a+ay�f.�������ͯ4O���,���廼��E0��3xa��8���N�R�Bu%��0�C�Nk? Ί|�]�O��2��@�:YQd�\:�0��Ug�?:,_�ӊ��\<�ӽE �&�(
	T�@�Y�^
�a�2�d��>��7�S��-^���J�4E� �z�X �e 9;����8��}�j�3����P)(&a�=iپU��Z`���< �)@L%�2�(�H7����q�,���M�}r+�� ���c�So���*S8A�ـ ���"�&ʛ��|?[c��]7K�][�:b�*"l~I�]�K�5F
>�(0'�$���I�����`g$�+�ٽd������	�g=���͵�l��{i�[ C�B�qi(�M5�����a�Q�.;���Lr3�BH�;�(�T�%�A ��Z'`��A�*0���8r�r����ecf�8ZE	�/�#� �;��҃&���������?پ����Ȳ��1�8�]b�2���MH��iz#Y���t�/��h�%F��U�1��f�Շ�\�Ec*P�3_J��A�y���`Pe�&��þ�O��@��8�ï,	�_T՝n�O�߉���)��O,s�	�����ڰ|T��ѡ���)ڭb����ej��G�b�����3��ե��G���d!j\�}�q�\�;�3 GT�~���%Rx�ҍ�E�<����ŷԍ/�}�+��d�<����f�$$H>����>/�H(������W�rk��К���_~T����'w���iD_�Xmϼ��\b��,נ��O�#%RC������,(�B�����%S��y�<L��L���u��Ge�g�J_��u��T�t2Snq��B�Mm�ۧRk�1>v�e.��F�9B�c���Rθ�H>.6�Vj�!E�"�==�>`"����$G�Ѧ�u��!�S1C���x����X�YRB�PHj�ڃ
����S��XoKE5g4b��$U��8KTПj�'֠_Y���H��׻��!cA���� ���n��5U!�02CJFIDn@�*�h�]/u{K����h�ԛ ]�kª�F.@�)d\�˗�� �K���1���Q0�\�$�(
j�l�"�)�/�kJk2xC�M)�O��t�&�p�u�&᫮��;N�l뼺�Z��r���Ȃd7���%�G�Qr>�VBU�:�ǠAuM�j��5��=�~{o.YS�@�����,��W�.�Z:ޥD�yP��V8�kN�����"۷��X�|"�^�r�rO�*���d�OҮ)�O"�~���z�O��Y�E��y�HI���E5�̱J�W+2�32��1���"�C&���>�c�قU@�B=�E s !�T�x����[W^􌴈ں�'��l폑<:5�i[��BX�!���D�b�O�3T�a��\�� ��٩��-+i�_~����>�c0=�Y53���=��vQ#��j6���������t�1�c:q�5�W�ųsؖkt��-ҹ�?�@�c(pX��9�� c�6�4�opD!L�+8V����_�0���3�
X��9�Zuŷ;������(@���%��B�l����E�5%���>���0�����&sqlA�tU�����E)y��o0���(�+Tv�X��Q����1�M�phKƿ�V�GV�����<� ���Z<94��)'���jlY�5'n������X;ԁ�aW��$�< �_�ԅ�X8�M�ٌ�y��ںC�B��w�C$f�s��[�����k�k��!���:z������V�����K��oT�(|\������{S9_�'�]w����q�����m=3�vh��V�����7S��0 ����=͔�J� �|L���.��Q�X��=L���n	#a����,2�ٯ�_+�F°	xQ�oG0b�
@aY�&�j�D�wl�
�Ws��1M9�n$	�b�[/�,�Ww��,���}S���L��2�m}���Ǝ�g �LOb%~y�8A�kφVx����� ~iR��y-3ܑ�0o����8��S�Cha+fǮ�-Z�3�/��� ���5�s���B�׶x˭���'����$�Q� ��թ��M�e�|�����E�$E� 0��Pe(σ$���2�����j-�&�{Hp#�J~轰K�a��3�@\�;�ӥ��f|��d��W��_/�	�p|�������mE���B�YF6BI��GT*�)���0�ˎΓn^���@�S�Ԃ�1Q���z�����������fz��*��$�|>�1��֨�����{v���BS��H��2�Ju�����g�4 �{�bhR/��vx��R٩�M�<E0�%H	Iɒ��↸��	�7��K�`s?�M
9� E��CE��V�%R�\�}�Mʤ�E�����xKRg��Rj�0���+�eԘ!aWEK��_��5u�}��8�H��W��	&0u�"�#^���V��O>#>��by<11�%�x)��Bt �~ %ʍ`�NI�O�B�w�MD�" &�9s���E:��B�]1��P�ȱ��o2MF�R��r	cn�eqh��cz[�O�jc����t���N+M,��ir���!�eK�S���SX���������]�"3
f�<0�n�Q����n�m�>���-��DO:]�0��L���\�$��M}y{1�HS��4�n�|�5R[h�n{���U3-,���@�#}jM��t1n��!��9�#[�G1���G����˄�5�ږ�R����g���T�)�"�����8��e��JY��I\bq#���:�ˮ��	l35��E!�?ʝ����jwjT0�Y����L���L�@c5�� �E޳�p>M42%7�[�xzg����7r�U&F��E���U��!�k-|�d[�t
��٠d.*	T|oR�����g���(���� O#ɩl�͊@'K���&H3��ɘl���2DZ�Ǐ*8l��Rӏ+	O`;�*Nq(��� �[~�|�R��uR���an�d!HyH+Յ��F�K�>mc����=]��d��@p���3OQ���Ay�����|Y��ۮQ�~u�p�������\��h1")�A��|\ȁ���R1�G����bH���bj�ȑOe/B�*��;�Vh1ݦ����Ye�;_<"
�I6�a:@�Y��8��?��\�8YU��EU����ck���H���.ؠ�}����*ֻ�)�3F�8�Jx�6=�{�.ϫ��ߚ��&7^%�B�xA.�3��n�l�i{��"�̅��.9N�� ��'�Z�d=[}
����V�\k
�?Z%-��}��M��Q�*�"<֡�H�	�lp�P*/���0�0ﾻ��Wo�����l�/D��� �Ӣ���e�ox����h���K
�"�%��NUB�n&�ӎbD*��j`��
7�E��mVZ�͍ɨ�1.�cd��[
�tb|���̭�_b�| w���P�±�͓��>CF��/� �+��H_z2����*��/�m/R}|KO��Y�;��dmb?�M,�s�7�zAK`�o�,���Oڍ]����8���4��醄ȹq��}N7z�;�_����A�����B���h$��u�������M��b��*��5�	Y=,ܥ�yE�O����sb�{Xkī���K�C8��p����SI-�41e`o4\�V~?�3�p���S�����5�	�i���H�����<�8F�.ݚ�拞p��N8e�Ѱ1㒇gU�S�8��@�żC�@��w�Ņ����/��-�ؾY�R&&�&>+PA&^�n*!�E�h�U�]��D2�'��ZP���<�j�n�3�X9��P�'ۯ�+�H���]���!�7;b?"}G�gX����s:��D�Z�Э���,B���qV����ҪO@�S��4��ET��6±�" my��LO��X4�y2��J*X��7!nq��T���uw�7��I
������ѝՊ�-�w��:�{<���{�AB�$ɖ��)n��/��ؚ��j�r�T�!BZ����3��N���;�L_���ÊN�EO��(U�9�n�6C��,U��:r��r�O���y<G��<����p�z�z\M��=[�w�0�K���*��N�4��h�>e_��+s�@�(����,�5^t�-��Z�V�^�.g�Û��]�O� �u�I�����o�#��tr^`��(+DhJ�q�^x��j ��X�:|��=�\�6x�H��Q�)���$�:T��W-ڮ&.{4
�3��ʃ���M����#-�םR�9L�ߟ����}]��إ�Q%��N����w��=e�y���{0��_2�f�����ȳ.r�Z��?\Ƴ�n����"�s�PSHV�N�h���3�z�<Y��@�(Y��%/-��N�M�F�G���T�8���*A�܄
�v𼲱��&rMr��#7���1�E+����NQ%&Ʒ�>].~(�~����� ;��C?����93҈\.Z���������\c�lu+�ٟTX�h�G�$�c$Q&����vI���`#�~�	�E���#<ڧ��v��q�Y���q� ��Q��Ɲ�����x]Ld�V��q�a'��^�Y)�4W(V���JHz]?ҵ�o����(��.��1Q���-̼����󘓨Q�gKx����j쒩��o[�����=�vO���S��S��w ���Y��]����[��e���.S��"㴟�$���m����H���9\9ph!��l�ί��b�����Q�'�~UG�|O����@����x��\��[7@����76hzT�Onm9����I�e<�G�O�qt��c�	������� ���
Ы�k�-��}���c�}���v�}wԗg<�u���}�	z��:Ӆ1�A*r�M�=�&^��z�{��\.T7sh�ŀ�U��0��M�x�O���o>�NSf��&&�!�nꙢ���^���o�3>,�'�i�p6>ax%�}|]Y]Xz���(����ty��D�9�Y��(-��3$9]�H�O���:�`�#�4���=�:dUa^K�@��j���F�͏Hأ�4x�~�^C�2�ʏ�<���lZ>֊��_!Y��}m�	��m��I�$Q�����`诇Z���N���R[uiWHH�C��og~m�]H��m�}���d}�n׷��Oc��w����~�.Fͻ�q�=�A���h�ϟhJ�g�A2���׾�l�5�/�*���ŉ��K�1�����+w�x��E�b����������0��S��ǂ�md��������L��L�V'|V_�2� ��M͛�~%����n��o̱�������T��nx��M��Aa~��R\%w���	�v8f�H�$�.6Z�5��㠂:��vZ2\ý��$�[�jfŗ^��3�	PF�;+}TÛ����dOfm���QЍ�P��_˄���E��ϸYP�$��qt��3 ��-F��_�'��e�8ShF��v��Qj��0v&��te�Y���)t��.�!���#����+���8�B��@�Xx����>D��d���H�!�rɏ<�۱q+���:v�����J�ŖY�rh�5lz�%ut^�b�Xqb�Y;��wᖔ�43[�q��U<J���hZ�\�Ͽ�+ �>�PY&|�X��Z!��dF�>�X�PnvP��<���,n� A�e�&A#F��Vn�ﯸhyD8Dgx�0��yybI�D�7�.]ވ����$�	K�c�"��F�a����01�v)����Ya���C�Ptfy��P�??�4|��Y^���:r��M<Eg
����mŸ�DSSS��!&:B���S���o���zˊ"�V���nA!��?����Մ�a�M$K�\|R���G�yҰ�z��N�X�~�P��X^])��.�PӇw��c���G���3<�?���~|�{�;���	 *dH�"�	Nn�VC�����-�7I�F��S���y����$z���X�\�#Y43Z_u���V�II��Z5ƻ;���ͧQQGv��_L���!�	�h��D2M\�ɛ4��Q��Jk�@I
��]�DO�E��ij�_d۸h��C�_��d0�ְ�b�>��O�ͫ\|�Gk�=t�3�#B�SH���I1(�^�[�D��%+<������Tc��̓U7���Sғ��`JI���� �ˮ��A,9�"�r���Fzg-z���'	��aᅥ!����Ѐ��N����^���έF��q�(�^s��D:�e��R�*G{(���xȍ�2������ �����IH�C�̹zrNY��.�f]]v���N��L!�L��wtI�@&%'/���:�)��o�y��Dm��[yW�9r�r{KXԠ1|jt��7��v� ��i
9ǭe��7�rql����	�\s$�Z��ֽfO�?�������ɖ|��?�̤#i�n�Td[(G��:.��h��$Hcd`)y���B�pXA�v�f�H��Bl�D����M��n<�o� 3���������~�r��7�U��`��<������C����@���AbW�,�'t��x��ȽFJm��b��T�k���l�<G�o|5�{ޛ�}h;��N(�1�y�I�>9����v:'�(�wd(�W��c���t�5��8�nJ�g�S��5�[�g�l!�Ą���Z����o!�\=��0���k6a��&��
�e�Ht���R��6�_��mSK�rN���UPa��oB�8�b�?�,>�T�z�\��f'/=c8�g��UP'*.�&ީF�V�y�lfļ�b�.�JQ���g��TǓ)p���,[@:�^�@F�!�|3H�h@�	%Ȭ�5���_!��B(U?/~2��ʱ�-�k�	��:3�J��kW2E���ڥi6�=�B����\E1��\Ű1���r�̈́���4;�;�"��6sd��k,̳̱���o�1�C.��~	>�EVQ1�~�}X�����W��>p��C��&��:U!ʫJ�U��.�|��Ј�Y��^�
b�Gz��sg�> [B�ZҎZ��J�;�V��ac��1Y��⇜<e���EQ�˗+6�T�	Ss���lk�u	*hp�$��Rru6�&U�A^��������rw3#Eȩ��g�X�qO�/	������I4\�>��g_B0깽c�*��e����t���C�<�<��۝B���S��c��N�s�xs� ��v�R�u���xb�mi ���5�ࠇ�p�c3��Bc��u�M�"��ŽZM���	�@B�F��5�6�0�@z��7�����{^�b}�Z.|{�t��4�4�쀜)8�4��q\��ċ+P��7�0��/����JÖ��K*V���N�R,�� 9�}u�ܪ��:�%VᛇgA�� m,R"�5Q���y�N�]�W��\hx��י�~�ǭ�C,t5�4����
��)��+�C6����`�c�e:c=�&��
LOi�|{E��5���чB�b�V��FU�^*����q^��ܗ�c�'u��u���m�Nl��s�.�X����pM9���I�q�=p�1LA���8�/ܕВɣ0�~Ô2���܆��Y8?>#��E���%ֹz����}l ���>x]�LU|w���$
c���Ae��D1	��B�0z���O7c���/4���j!=ɓa�hc�I����&���b��/5͛r�m��$�pR/W�?+��/�WW*�_�wZ����S{E`
Ի&#K|��ر�R�$@X����E1�F��o��\����!���;g��XY�HLX`0������c�;���Y��l՚�.�)doڬW`L��Ab)A�F��l�^ѭI��o�UF�>�9r��A}�؜G�}9���D�n�4����l�*?h�Y6�z�J���%')����j{ &ξ����#j�i9���%��o��sii�R��:��<$�n~�������_n4��ƞ�B$��;���kl
;�4��{褅�X�.����?Y$1�[tN�b��h������=�E%���9bhoLK�,:��������t��V�Ƙ��?G�{R�6K��'�2���f.�q~|�m/ױ��S �8?JA��P��q�}�vJ����a筚趘���+E�x����tvb!Ps30�Ÿ,9��!��hD�e�%6�GW�����$�L2q��?[6����yI��XT�዁*[t��9v�۾�(*䆧�&��ѳ�>|��sИ��ֲ�Ǩ�<���e[Q��b4�y-��5��
��G���zwO�tq�s*���1^�g�fWL*(�M���̱m�e��j6�\��4s�+7f��D:�u��������$2)ה��;skh�&@=�!��g1	P?�!V�{ �A�D�x�2��ﵲ
v�e�~��f� �\�@��zS�����
(�)��8a/��c$�M��`=p� I��bRm�Q�dL�� �;�I��O��e�
��R�}uZu)����+�B6,[��R��Pu��(/+5�H��K�����1�U<��:$�}�[��@�ҧZ5~���/;�d&�t�z�z�ӡ>|W��{a?�
،���`�-f�9�c{Ln��ɮ���n>
b�.Dѣ@�+�weDG�&���6���Ii�%�[�����ʻ��c8��CqL����r� 
�`�vy``�+V�� �D�t�9�a�{e�yXF�TQ��+��
�)Q��
��F���Ћ?=j�
8o�)��܌�|���OH�^��03���Z����Bg�塄y��E�s5Ǥ���:�V�P6Ķ�݄�H3���r�4�nxde�En�Ք�]F�d��y"�z䉣n�%Ć�9U�	��7�";����؍z'���spdf�#�;����hZτ��>}����
[i*�����ZI�ߖ,����u��b�A'A���Ao�>E��)�r�&GVG4�#�y�&lA�ȅY|�@Δ1�\�~���I���yo���X3]�[��d��(_X���B:��L�	�2[��{)�*t��ŭ-{#��d�N����{Z˛�Φ:�P6�����~�x��˃�컡���MB�B���i?��@��-�d�ݴ ��&�ݖ�t�6�q���W�;�{�ʯh��M�<�ËY6B<G�wg�0�RU�f��1��T��5��ߛ�:��X�[�,�_߶�z�]Ew���}��.2����jУ�A
��+��� �3�@�~B�Rk��WL�r$=Y���)x�>����R��@J5	���0�%+��
Ufu/��GKF�	�itZ�IJ�����{����/Y��Uot��L ��~8o�ūVx�HXK��'V`�ؚ��"���Xۇ�,V"����/I� ��KK����&�P"�����e1ݝ�r�=�ےMuN���hۮK}{+S4i���s���/(�%9L� }�v>ev����[f}x�� ��n���q�.�2�ۧd��{��yl$Boi9,i(�P�T�p��	R��\,k-��t�~#�@���#�Z������N�,�xթ�nkk�63�]*׉O���&W�KPps�(K��B�@�9��CSy��� ����p��l�����`�������V��g�jS�5*JȊb�!.����跙8�]���Bp>R[͈���rO��6��K����������Y��*p��.�6����2�98�M�(�%ư1{���\�9�!�x�_�LV�.v��9t��2<������Tx+�#�����U�WmC��i��#��L�p����׺Jϋfl�,���f�K)/�XT2�9�5��ñ��BX��&�A�m��j��Lq�M�{kr�fv����7�!U�Ӄt�IO5~��[4�?b��E�;ҹM����qR�.�@�C ��R�աr��&���Ȍ�Q�q�ެ��z|h��d��b��!M�_�x���!�th;�4��"���cfJ���Ҹ�x�4�x�Ug�N0
t�/�A=�'�柹��.E6@T�/ھ�^a�|�˼2�2q���JƽѠ�Yb2���S�_g�=l]� �	�!�J!�l��Ϊ����KS|��;V� ���*�cr�X�����d}O5��x?W��(�
\7��� �)be%h%O)O���B�bd"���C��q��4�=�����5P�EN�S�Ă�l%c��K@�A��&�� �MQrڮ`�=��t�i"II��U�<�y�D�%��Ϡ�+�����5�V���هm��0�%^�G��C�ҧ\i�3�*f��CTB�ث�c��慔��fk1�U��)4�6:��;�s�����=�M�>�(�$$����w��`2vX|v��n��)�	��]:�x8�]G��������f<�?U	0����4$����2ʂ4L�C�$<�C('0����R*�Ɩ3�Rf�O������)�/��!����& ��7}D�^�/�Y<�"K����	���o�_�����݇�Q�])����ZH2��w������5��%��������gt��N#���@[	����W49Ҙ���Q��HD�8����x���o��萯��tb�?3!�|��ɞS�m�r�O���󄕯�su�t䥐��q$�Z�sw��9�g�A�j�1;_���9��+��c�N�����'���5�]9��{J���fD.� �ͭN�������U٘�R�z���#�]�.�\�:�~l�P|��#G ���}5��є2�<#_~}<k�}�';�����o}���������{�[��:T�#`�Y'`�P�LbD6!�LU����?v�W�x	��;�����a�9�^�~���d��]��4��8pl#vj��.�C&<:��w,943��&T�����)�/�1��W)\ ��"��FhR��^~W���G�����ҎS��Wƀ)Op���W`,xf�hTs�{-w�@��M9KA���D2YO�K����5˿nν�������O��n9f^�w/�?��7Ҫ���q�^��&�%z�����P��㿨�>礼%h���?��e�?�i��Dޔ?�,{Zg(��X�\���Od�|���=VW}��3��AD{6MY���E��l��ej�I������_qt�q���� I�ѽ��b���7r�4L����r����K^��۠k2(���M=2����R𫧖���lx=� ,��ĝu��{Q�����T�Ip'B$h���h<<�n}f��}q���y������	���~�*1y���&'.H���e���Z�̞��-�O<ʹ��ǰ&�ƕ�;ɡ�zg��V�΋E/hӚHy�;`H�7	�6G�/�d���hW5�o��sLڲ$ ��/� �r�̵6�{ڜi;�Q�m:��|A�ȅ+w�6�mTx�����E��7 �r>A̾AJe��,wJ��C�[7G�oB5bp1��{Y�#�B3�~UϽ�&�f�{����c�-����s�g(�����ŀ���T�YE�m&r�%k @b���b=�JE�o�l�c�(�!w��~�3�6,�r凴/��{���ԍ��8.�|U����|�ZV�D���`��3� "6�bQ��ko�� \���c� @)VJ��\.תQki���"�vD��- 3��m�$�!���@s��tK�5�%< ��A�	Ue����$&�9�OG1����%J�3���w����S��K�)����@}NA��z�Y���8.�J�)���2�(�'�:�j�"C�/v�vջ�`��Rˠ�3���]�
��q�%?%֞��,UY��j�VX�s�XK��̑��``P���_�R�~{ۅ�X�g�}�a[�y ��=V�0%���z�GN��F��cwj���?���B1��h�"(�6�}���V�������ŖO�kSNE#E���X�0O'T�A��?�-C#��W9�c�"h�n.U�����8ҙP
�	��.i"�*�c}�/2�Dz��=D��0/P52��-ߡ�J�0:ێW���*ނ��nc��5���@w�Cۆ,'AA�ϸ>Ĵk�9%�ަ��'���^Rt���E�v�ιl������B2��N3+z|��o` �*�y�!)��2=�$�y�&#����"e���ב�?�P�%�ΨY��� �^�<�Q����e=E6o�s���e�m*ܸF��F�Cpf��r�{�Xl��T�;Yq^y��L��.��إ>��-���mP���2�3V�M�O6i[�21��,.f"�۩(Yˠ/0��.�����o(�L+������]pRJ����reQU��~�rO�-�V�󙟌~(\��bp���A�a��%jև�(���;��&�����n<;8�&��H�j0�$�Ռ%H��.H{B0�ͮ��µXKQɯ�+]فCh�U���}p�+dj��t0ӵ����ZT����jS�����R���x��"���ʨ���ό�,���&���sQ��T�cP�n�Eڨ�}`�@2���O�����^��tZ�x�!uo��g	8�K�}�v��ARwY�v!.�by���/��վB7���)����9{DZ=w%��9��-�͞�E
� +�?����#�w���V0<�cpX���p5i�o�vkݧZ��М�߮����H�)��O�R
H0@5A�}S��Qoؖ��Q.���85�qxU�m�:#?����Y���^�$��9�P��;:g��/Qy��~�n�5��^��i�����hS���?��w����J��nW�E�UgU4󞄬Uyͼ�Y�8t����� �};�*'�QR��w�`Z\٩�JIWSg�̿�`�}Tf_��6?e�t��t	�2�ɋ���3��oI�w�b�`��!�m�2��,oJ!��4�ڧ����K^\� �9IZR�o�e�s�7�_�ڢ��%��x��w!f�47XuL��c�ɒ�N����Ҁ_
��R5"���Z�(#����?��D����BlL�(�9/�5s�z�i����j���֮{z1�����6�)�,,wAᘒ�p�C�&]ϒq[��%�盖%3���k�b����=<4kz���+F�$g
��v~��R��k=�tE��~�|���u��.�C_�-��������m�*r?4�W�#6�,�U�v�xv����I�7��RM)Eh~M�e6<z��ց����
���Nt,�2S�$��/��9�j-�`p�.E%��0���:�X��# 
�=3:��*�����&ǃ��f���t"�Xm��׳��wM�+��[ŵ�pT��wv#_��h����t!\0>�C�j6W���`F��=R�|�F��MBk����oj
"$�3ӿ�5Ȉ��]�_�5�$"�D:5n�H���yz��d��,]�cHF�����ݷq������b��"ݱv��3]��к�%��c=����V��[�\(8�+�{�~��N��&VW3<r�7��fU�;Um�h��Ro�@��^�i4��U��e��`o�2=,a8����(��׀1|�)eLV�����w�]����7<�o4D���K�����v�t�9 �"����׀*�f�t�At��L�dF'/2�8{��C�:G�������qV�o%��s0w�R�������r�Ur)WZ�J��ap�F����c��~�~���疚�>cWs������Au��\����ȋ̸R��0G�U9^E8�h�s��ϸ��׆���|�li�����em1!�]��9�ܓݢv����c0��kΰ��}���٫ӌی���X���}��̞���wj:tt�_���O|݇֡�A��W#���" ��:��Q`RɆ���Ϗ� ���,�v���T�X���e5��tK�fJ}�E�� ~x�b0P1�Ī��2���&�Mg��`t�����?F�V�J���F��f��Aaţ�;=�R`�V�. Q�� 7O�뼎m�hRr��U�.��K���"��0E� C�NǓ�֊���7�M�K�u"�_)�=%y�9��݃��S}�E��>k����O���/��HĠ�7C�)����>
ןm�B?�y����C�qa��t��rYYu薳��ޭX�Qd��m5��ɮ�E2%��@{@�F���b��Ƥ�a�6��U�~�g'j{Q4��[��L7$��ZJ�Ǖ��S(�m��N >��Ͱ��,��٢+Z��g�r���e�I�*�]mk݂�Z'z7�ϭ�"�o�s��x�`5�=��Q�ҳ=�Z;�H�x���2��=���AV���<e����;���W�� ��f��eA�maa��(Z�S�mJ�*�,w��3r��O�1�'XIζ�s+:3�<��؅�d�V[��rc��`����z��T2�Sx��^��/�a����D�j�?�G�q)�W��z&��l�>����6mE�"�
�0�h�l(�5l�	����
%�{H�)�\k�w��ӣDƛƉ��<���"��@n�:^ZUR!���G�����N��92>t��쏄�!\�)r��.������V�T(�.ec�Z)��N_�s#� һ5��中
u��#���6��Y���[�� �;Qϳ�XܬK�B�1�;�ĝˊ&��jAT�|���	�C�X�6���s�IR�FhdZ\Ak��gO#v�&5���᥿==�C�j.:.%ш��l�AJ���O�(Ҁ���Z �M8��^�b�����#J)3}�>�C���P��Z>���8b�}�6�Pr�v��^�����bH�t�8o�U���iӱTt����[�Dao���o�T��"KO�j��x�o�14��1^V�j�KeӼ�P������`,�*�J\�U����i���b�$���V�Y��w��Tf��2���F��c���k��������R���C�r�A̱��,c�_l�=���H��4o��t����I� �!tG��i��������@����-��n
��ѷIK��,��T��Yo]���epף+�� ��柦���=��+z]��M��4]I�}i�����fɃ��&D=��+(��CR��c�\��J�e_zz*#]����q�ŉ#��YT��� c��w�%���R��5����꟫�"��;���#Gs��#�b�,K�)�� ٝS� �[�F/�Ɓv��@��ܟxk!Zc�[nt��5�pF���"�[M`�s7�(�V�\0Xh՝*�� I毕\�ߥ^��Ʊ,��h F��|�V-MÂ������3:. 
�hCn���f�e�~���б<p��w�P ��ǧԱ|7��kI���m?5��4|��n~#&gc6� RJ3��E�{Q�[d�O�4GV��P6AC1 ����C%��Rq��X��de��=����� �
s(P�׀Ȍ J�|��{�r 4s�#��k�_����@3�J%��$�_a�B�)��o�Tw��d�D$���WTw�4�%
	ic�=�T?$ߘc�HE ��*����(���Z��@�, ���&l��FHܴ����5cu\���)�^�%��~��2c���N)�q�E'�u�������MQ������ϱ����U�YSK�6����[\�U����w��C���cW�]X���8����?vK�}�	�J@�h�����+u���O�{��\]�a9��L��{�v�{�dJ�BT͏jN�$ٌ����D�6���F�;2u�����P�:��/_"*�h��Vm��pB�MH�i��Zlsv������̥S���.q粍����{\�Е���
��G�NS�ڜ6�"�)���_�~;�f!�a��+1�-�$%�-��k�}�sGK���0F�4�T�m����К�]{�O���x" �0�k��E;_���Ѷ�|�=�aW T���a�_7�zK�6�&�8�5�<<���7���a�أ��&,�YY�$/�"��7�ˠ��M�z �`�NJJ��%{���������t��x~ض��W{# �m<���͑s)�l��t��H��UvM�G����G�u��5GS�zϚD j���ρ*j�j[�G�]���y�����4G�]����NS	���������8�� �P��Ѫq�2����O��x�)K�G��(2Ӛ�!����ƺחY@&�G޺���?�)0V����eD2
�IY�%ШZ;��=Z�i��4�5���a�68��=��6�^��?��B�H�E�w)L���S_Q�N�!:��[�~�|o�d�.t��S�~�}���uUH7�	�j�:��z����k4����~Ѿ�6Z����*�i�9BK���eE�I��c
1n���(����=E��$,�dtO���}�l�E��:P�Ȉ��ON���c@�I��ar�Z���U$��$�3��6�Eoq���㪜y�A�`�CYP'�t�0��[�>����j�3���6��������� |d$F�%���R����I^�tG��^������2v�ޏ�'�:ze{�(V�ܬS9+u�R2��8yM��ĉ��h���Ń����M�s̲A��냲��PN8Ag�2���ā��$��o{X����&x�����I7�����72zX��A�ݝ��bϢp�`X���e�����Y�G!t#dֺD�-�\��<J�)�[R&��<�ns��Z2	��,�\Ш} œ��SP)�})rt�FֱW>$��ƾ�c�����2���
�λ� K��t�w���J���;+F��n7�,6V���.+Ɉ�붣mu�3Y(�6;&Έh��PKI5�A������x .��մ��p�1-��Mb3�R�lթ%m֌�гO|`�7��|�\�3ɚ���I�;c��I���u����2�����e�Du@m
 ��t��,�Q���bz�*(���
�6ڧe�S�R��[�w��Ap5w�s�<�  �
�,�^
b\����4���zLW�Tyv��3��� "1f��`ǚA�d�\Ѳ�Nٗ)֑L�7��T��[��E���#ź�:��:��n�+FK���l�c�,������ãY4������Ly�>:��"+�Ѥ����`2�c$:֣����)7��g���%�&g�.��.Ma�x���T:��P�PQ91�]���7�C�vER��J����NB4�VP�7�k�Y &��EyL�:��n	T l3C�b�A��	"3��	u|���s�c|�jB�����XD��~W��5���(3���D�2�R��b��Nl���J�m ���W��Y��o���i���Nof{���8:)�@ˍ��䪠��B��H�٘�"�|{��2USu����A
H���Q�2h�&ş�ig2������Gt��k�<V�KBh�c�����{,
~zִK���Y����}>�=��7�g�oB�#闏uږNػ�-�
^�ѡ��Iv8�2-��aPQ�S�0�{�R5l��o��.^`��tA��:"n{��(=}[���*�����c#�K��KH�tY�)��%B,���x4����p�3x�)��p����]���B�� �~�lc�c�э92d-*{�NT��i�R����f�����5�wۍm�L���L�*uk5�:�|�5��?aᬢ}x��u6�"�Y��1 ��ŖPxm��g[.��mM#6eo�7���v�O���W6L@��{��l�x�C��&J�f�'q.�κ1rv�嵴�Ĺ�{2��!/��T�<$�O�}�p�л+�2�A�4T��x:W�jQ͂g<醆��Qg�1<wy�gPg̔,n���k穝d@ΚƓ2S��j�����>��g�F}�	ʥ'�$7vv�������N��9g;�M'�ў�����ّT$�^����&��[��,�Є1T���C�{��Td��o"��Pi����b�\�4�a�BjR�Y�M��ڣxh��Y��e��A�G)Jӑz�fߣ��b`��&�h���Χ`����-�4e����zY�"km��%�p��R��H�>|5�w: lR,y�H��e�]E2�MC:��n#jB*����\��求�@B9D-oL���Q��G}J��2��3�u�%Z����9���
U��>%NQ�M��%0�u��y¸��q�Jty������3i�r�GZ�v��r�P�[�^�:����P8
cJij��\8R\�Qi&A����l�t�_@�ks�D�����OsL�~�]F�ç��*�m�c���!����ػ��Q
B^#����h9�|V#�� C�ԑ����:��1U��B<G���l�Զ-�̩_����i@�E_l�3�pI���s�kC��x�Փ�7^$��Q@V����@P�5�ﷆ�b&)����˶;a'���cF7hHR�1�"d	w�RZ��x�H��33M����cp�G���]��J�Y�^z�{�v��N�6`��2C�>�\e�.U-�L�{� GR|1�����p�Zty�/_-��Y�3�0�fpy͘� {��b���xhZ�Q�2������A�鑊τ��Ʒr��$��zUG!�7�bI{M�%*��^|��п�)4��E�.E�$:�W��x��K�^g=��4.�/&�b򺘌��d[��Bʕ�$_ 1↩;� o��Z�M���Pw��ꇳ�RPF�[�E�*l34^���H�H+��`���!�d�z��IC�b��\Luq�0�y=l�P�kӮ��ę`Z,(�gSe����Z*���!�NA�='��bNAl ���/����\������J�����Zwt).w� ���k��GV�Ϛ	��i��FS���/."d����WL�6�s`��Ъ�NB���q���d�� �Q���B;��M댐�&�
����Y�
�]�o��"�$���*���K��8���5d�8.C����)��6��1���V�E�R^��"�9Y��^=�>{!�a$�VyYm^�r��	9�rCؙ��Ea�.��ͨ2#[j�`ȨH�/I���p�pQ����
T;F`O8w%��Oy/r�A��Q�tϜ�D�A\=J�jc�R'�_��F���}�B� ��\<���&f���"oZ�}�����N�$E2����j$�GJ�A]��nm�k�
�vRJ2�$�W�l}�԰ߟn^��}	W�+�/�?���`ޣ�i�9I�Bo��+=C����}#2����́��?˖l��"����j�#����OJ�,.��«�f���R$�u�@�_����O�3��0�3��{)��Q1��{E}$V���|����G����<X0��_���ÍR�������mj{f�e	����K?\��xd��6 �`3�!>�yMaϑ/*9B;�h�E�`8���Ü�v����gE7�b�o����
ɣ���Fc]��1�P}�R(�5��n�h�*�H��.�=�I��!���?����
��Kb�D���*���L@W��kU�u@:�&;�.��4U
V�t�KZu4-ʚp���.Ȟ�0&œ�0w�A
dޑ�UG���>"�*ǰH�q{����{���Ev��7�cӢAq��T����c�S��R|	�	�d�lRI���`��ѳn�T�ʃ��)���Q\@�aT�� J
O �t��+��\�ԙ��$'ϋ�_OK��\�C��J;���|��Ab
�OFs�ܦU���a����z�
�R�]،C5���%�W2fμ����Üw�*�)}i���w���珁#�|d� ԟ먢���I��OI��S?:�ʃ��Q��Q���R`��	�E�9�kPJ��Wē�m���z�rK76�@tڗ�if	"�OA�p	����PgJ�ؚxI0�h6P�p��o���C1m�+�_av��|��+�xv�l[��,3�e����:�3N��C=�e���j)�/�I�����D"O9�K�;<)E��e��##�s\��My#�5܉�2z��Sè�
�˯d"�䑺x��z�i�qH�_d<R�7�C���d��c�K|��������U�-4�C��bx���&���
��!"j5����*O���,�����ů3�h/{�Oÿ���K����o7nHhHyv���$����0<��yQx�&��[%����uu�v��:�8�1�);���<!�K7:�x�k�8�R.-��ȏDF��1}�y���>M8*��-�o�
wU�*�Y����8D�=��T�.=�D"_V��_����ǳ����O����lvusܕg6���+37g���@y�� �S�mvi��8kH2��]c�v!����P�3���t>��	�G���DA] W���C�sc3�]���B�,(d=a!45�4_D3��~�'z�LX�d(�i7�f�<��|�������_ j��w�T�	�pq-���^�֐�Axo��د��#&z�����[�!q�FE@����Q��rlY_|ƒI��Q�2��T���
�ȑ%���'��J�U<{�~��
V���,CW��V{wJ�h%����� ^�R�<bApX'��SFV,�H[�L��'��&�/oy<�HA�#8�OO��J����k4�.�m��QUN�qV�s3��Q��r���6py7�Ʋ��/��ȞV��/.7��,jd���3X�z�_�"���lj���]ޏr�L�:��l�V1�FQ�J�i`q�&��mb:����|���k�Q�3�k��njZ\�!�L�e�# (!������+j��^�9�W����?�\0��9D(FJ@PE*rm���3��\��T�AH�d��.&,屈�U.\���[r�%�����r7�t�}
k�\6%˫����Y�'h¢�E&�~��	���=������4�9A�jw_���͍�z����i{�0�&�������^5��v%������3�-l0P�l��Аi���FfT��X��v�B����UJ��`���B���J1B3ILu20��#�.k�i���Yi�Q��v�mֈb<{kD�z������ZZ�rK�]����ĺ��g�~V�u."s ��d�~6|�_�vH��|�ԒЄh�i���m����l��ڙ8���!p�H˸���1����&��@����&;��9�����׭����vE��^�7 ]���m#���fe��|��b�wԀ|�ٔQ��o2���hh��ްu�9�< �%esipJ�l�6�QJ2V�:?��[qOH�ԍ�Py��K 85�Xz!q\E��uX j�=��7��['�UF���YxU�o�kP��!SUC���(4o��w�J��hƬkbP�t _"��,:ɍ��g!�)g��q��[�%#(���
�	��Mϼƫh�����P5�W+I5n�v�;�E�-kD�/�4�(/�sA�-����,� �FAF��Ap�j�9�u��E6$������*���OW8#Uf���ʄ����=Ml���Y�r�m��	�oG%"II$��?Ś
%BF?�ђ�o%�ߨ�͋ ����E(
�ᯫ���=�I������Ω*��|)��Ɓ,u�[p��d��c��:jAH�J�H'|.iI*���."d?�Bt=��p�Y��g]ve��lz~²O@�^���<��r8���D�/�2��m0�fbj�85������R��+��������4&x���3���+��?,�|jE��X,��ika��1��V?�Ե��V��J���|e�&��t�n, �p�dg>�և�MOs��������Rg�\�d��7��!�]��߰��~�u��E��F�^��0R�*n`)B�x`�*kݞ�����(<n� ![q+?�%X����n��NHU��&`q:dv�k*ۛR��0f�w�ҕ���Gj\ܒ˅L�y���7p� U/����O��b��Pݽ����M��򫹸H^��aH;���;3Z͜�O`���OpTL�~�*D��8���z&{�S��d�0�����<)`dC�~&�������1!�������:����]����[��<~c��
�Լ^�t2�*~�,߱m�W�E� ,Dr���:�Bj-���	��#�T��I���+a2j�����;4J��?����4�t��yb�2�l����:�+ÙC� W��L�@��S�����;�#�]��q��B�%�`���
���,zst���<y�;�����KFT?���j�ۓ̺"xק�f]L�İy�t-M�q.8L%>�W���a���*y�����c2�l�ab��,=w<#혫��F<7�]�KL�i^�Z���f{��㜵3@��b��EUIw
s-99��Y!�!�R����3���5Q;C�ށuɷ�7P*�PMlzc�h�3F��~�(��H}�d�E��h���o����ڶ���f�a�Y�NL�G⹘��(�գLq�v��������./G��/�=Pb�}��6����6-ϙmk��5
��D"��{�SO�~���vu����4Z7C��7"8�{A�9n�����Yt�NLr��x#�oLP�F�k����nЃ��
��_]�}ٕ���}�dY_N��jA��W[R;Y:-�����u��_�5�PC,���h�c��	"ꭝ���l�V�+���U����/����e7N�Pb���T�,ՄoX61<O����x˜��l���=>�	����|{�tU��*�`g)�Ĥ�0)E]qߟ�*C�zx5<NB���9���0P1����8�f��|A��Om]&nw���<B�C'丮S��{�3wѿ ���18T�%�' |�#:\Q�	,Ǔ��Tv�xn_T	�nr��'��@�V��5;|�e
W��X�Q��I�g��g���M5!N���q숱22�k�#%��_�Q�8�3!}1�͌�@n\�{��}��=�$jk����Q��m(�%�려��Gj.�;�Al�I��m��;�rM�w��{S1NJY����U��5��ب�W��pYj��0�@ե�M�2�?�ۛ�	|�SK�A�M����n���ڧv؄W�0�vm8�f�A(��p�WR�"\�f��֋�����*sv�Rc.��΍�e^C|%T#o�#�3r�����=����,'2�:�Vx�TÆ��	m�8��#�!�d' *��-��UCS�	�j���5�^3������	�CׁmsH�>0 ��]���=�pw>�L���l^ �RS��G�H$�4�+i�L,�^��n���{�Ή�Sg@�;f�����/��
����N������D�~z���y��rEgr�[mX�F�x��)ѓ�<����U���B;Ex2�KA���=,A�ȩ��-xG�_��m���Td��_1�^gͨt��ɔp=��!3��t��U�~��r�A�.����]�&ku5lq��3L��ȃ���f�} ��
������Z���&��a҉ `��G�}c�G1����l�.��W���L�!ȫ���s\jz��2hB>�L���%S��%j�6�l���ɚS�?G�OY�^�d8.� ��؉�K+Rk�����v��A� !3ڗ)s���Ph +�(���q��P��Yٟ��SmT>`^I[�1)M�{*V�{�8��B�{�A��Ҳ�6d�����,�i�{�uJ����=����K�À�p�0�9g���ڵ:F9dyu�}��r���RtEi���1�v>d�����ZL꒧�K���'n�Y�L�N۔.)��!���4Jqi'k�ٮl ^fr�n.e�������������.7��i�W�|d�r�PfoѢo�P��zCK�d��}E�C���K��;lx�>2�������du!��ck1�<����
I����O�a�h�Z/�l|q%Ϗ�%Jr�R�i��43�;X�&J, m��&^w��q^'M}�h��ݪ�s���ȊЦ�aZ�e�4�l<��/@�<�����<Pߠ"����K�\��坣��䓭\�/Z�K)MZ������:���֟J��J���ݙ_������f��wlx��L��\��Z�Ua!�1/���~��v0	T2��h fdSlPB�M�MmtkW�\�]+?��r tz'���2mE��f_oq���C>]��t��"�xF>(��Y,��VW!n���I���mv5�l7���, h[N�<�N���b㰛��P]e+:a��k�4x�tB�џ��xs������DC�4F��?��+��A�o#P�����O�z�j��t�ʺ��x�G�b�M�h��u��b��IS��2�LL���n;�x"q2��������������Kvq�;I(�W��P�W��Q5%�^��x�_��ܝĵ����t�ߒ�^�֢.��c���ѲԪ�-��p%�-\8d���B<f7$	�\��jR���+mݯK���M^Zg_n���L�������^a��(+h�_|�VFpj> N���),Om. L,��K���r�m��Ѭl�& ,ށe�5��9�r ���~a$`�3=GSMv��iA�;��Q:U��~�*��߅I�D��B;pDcQ�ڷ	�`�񊻼H���ε0(�ć��4mdB�����M�Ńˣ)��v'e2ӕ`~Q�W����ٲgd>�	��>��d��&C_�F��cb��A�ơ�$����q3�$�:N��l ���L�b��A]�����N�%���_*}��Dӱb��M��"@vj�u�R�G��b�U5nb��`��rW�@;�ˠ��h�q���g�<Cdf"��P���Y�ܺ���vxi���$�����F'��%��@������*Z1���<�y��L��r���~���8<[��\����?�,>B<�l�"�C�C��f��YOM��w �M�$��W���i�4!3ߌڣp�^4�:�!�{����rfx#�����GJ�O���h�V�ub���}��V£[lM�1�?n@Z=�����2=��11}�	�L�{���,.]��+�����]y����T��� Ul���#u���)3���	�l���ًR~������/�����#�wX �>�D�d\u�{<��=�A�Jdv*V�'���C��u�]�g��W�[�[�L2I�A�����#�W��1%�ܡUji�KT�����-i���*7��w]�A���h�m�ȰH	�CA��!\H<�$c���E��+K�E���F�H%��>��P�5I�%&$��T�(;U���I�����J�T?_�~�1���d.�X�����%ok�����n��dG�M�#�Zg��N�n��q�nް������!������}*�/�2��z���?�>{��}�U�\3���@��E�JN�Al҂t�p��ufߩ��-�wF���>�2��=���2�/��u�b�3X�#�_J�[a hʺw�4�ͮ��eDD��k�*����m��M�jW���P��)�I^���1n��SI1ﺅqL��:�}+k��mi1���-�fl�#�W�Z,��<�ങ/�`7`~�'�f���+��ݜ7X~Oe���w���`�'.~_L�s����r��U���c�=Z�.R�^����C&�<B�[�ozO����P��aOW�9�~,^��"���m�����qe-<�����fKĔ���jN��C����G]TZd�c�e�Z��6r��Ye�N+�wXw����Eް�]$TD[wp����pA!�KP�4�^���π1O+��hg��T�PxA_-\��8]����e��[T�v���b�U�e��J?�;YM�w�
Tm�k��m���x1�!�x<Z{4ET�v�q1��ܤx<YD[]O.cdCB<�O��k"9������������Ǻ,?���i;b=���ߕ�tچy)��i&�_��҇���g�;�n�D��l�Fm	E�w�.۸��I��3"9u�w�'�4�&k��;8Nkt��BB��;W��b�,)Y~W-A9ײ�d[��. *��LX�u��m�\��Ѝ��� �Ö�
p��A�����K��w}�O	��K	&���o�(���=��-����ɗ��g�		8~/V%� o܊�����ڨ��Ŷ�ZVT62��|82\(���X�NX��*rQG�/Ӫ���ĠuD�m�?�� J`��s>\���G߶F��1�3��av+�5�[�b���4�b�Ċ�/�n�5�Ҥ���R��2�ƺ;I0[\�ǟ=��3�
4ͯ��pKg�D��k^@�t��"� x�cKb�87�Ϥ,o�jw$1@�{�&����� ���\�����	��کB�yIȾ��U�^�,�P��X�&w	l���( n_���*�͵)�� ��Ykq�i�� �6��D'��@+�� ٭����51zBB�B<�m�c/V'�ok.0�-\ S���ǲ�3D-��2��舦3��+t%�ȉPr�c��"�U��l���A���������w�~l%-�nP�[�2z���)�
qߪ��A���P�ʔ-���L�u��o���78CN2��XW�!�{k,j��r��@'O�;��Y��z%n
{i-'�MN1�(yf��F�N�վ��QM�m=͞Z���F��l9�����-��n��PSN�ח}!sV�3�h��C�����i���F�2ו9�a��\��@���" �u�}@�b@�/X�K2��q�!������{x/ۊ��)�1�h���_��+��4d��C�˒v�0TAG��� {	��L^�뜢�Q�a�8���Li�����������9�����% �9�k@��M�߅��9���k���8��2y�2E�%�ڒ�����sr�YB�Z��.T�\���������^�[��y�G��j^�Ҝ����M��T �����K� Yu�T��`��yr&��r���R�]N�[c7�j�4T��T{��k8΁ɜ�[�Z�=���N>%8QQ�ͩ�o1�����[pF;�����8(=�J4ŉ�9��A�R����#�q�5{&�u��(�W"��?�VRO�fE�]/X6^�XO^��rww���~jlz��ğ��*�%���ʭbӑ7	y78���@Kvrb�B���}�$�a2���[�w��V���偐,R�j�
{�MH�EЙ���lx��G	"���A%�=�#R̚8���	�w#�c� ce��5���eX�(^h�H��g��ƈp���G-T� ���W��*�E ij�18��>6el�o�œ�x3e
XZ�!�Pȝ�ʎ��㒺���[?"ZY|�h��� �u��D��H
|(
T�j}h���F�$�ޓig���rI��6���vs�{�9Fa�X� Dg	�b@�\頻?[��0�U-_���ͣC��ʭcM�"6��=|����m��M����)�vEq�ve[4Cv���|uO)@5�Ò���n�&wa�?ߛ�إtѫ� ��_C�3�o�g���Y�(�4��I<�9�@����z���N���fT�,}�lX���N�=�Iߩ��_R��DӉe��!S���¯Z\��0	kzc���$?tw+D���'�۫�/���\��,��g�d*��荹۸�z���7����W�,d�oR����0�# n75O�x�?��' T�n��+�d����vpOեf��g�HE���7�%E����Ǽ��]�XF|��e�lIgjf��$���Ɨ
{��<�"���'77%�E��8dqd�`�I��¦D�<f�����`�_]�*�t8��l"^��'�q]8�7�'�;\	�����Z���P��/���n��E(:���
8����Q�6o�&�>7�-�&:z:�Ӑ�6�&��-�Q�X�_�o5SfI
%	�
��  _�.1$��1�san�?�&���.e�k�
v�������k�A9�[t1�Ub���oW�K�ZuHw�w���3(5C�e�z���׺�2{�P=�c2ixj�-)�ӹ93��c!m��t6�ﭱ\��q�0��OX>}S|)�ٚc��e֙Tu�Kl�H$�NT�����.-ܶ��$8��{`Jt�6H�ܟ� ������O��B�%�0�sv��h_��^%آ�D�!�@��T���4p(��	~�jN]z��*ز\������C��fq��4�Q�v��9A��eߑ��71	'Ix����w���3��jD�M� ~ҳ��� +�{�`)�)j�A�VDM���g���,��}{�A�c��}J�	�,�dG�g�^>�`^�lm����C4=���˧#+ �:����5��]�#��eS��Н�d��N]�c@o����|�p?���������#��y[,�e�/���d9��©7�;��E�Jz���rd�
|�[$��rD$5�~K-�+�[��U�+����K�" �k����%\�,qZ50��-�ҁ�R��F�d�
�J�`}��U�W��̈́���7疕jML^�%w��CДwˊ�TR�VC�9{�K�ܲ�R��R0Z˒;|gM�5̵]W)A�k�{�];�����UѫN�TCT�����n-��A�=��zZ�e�@i̝��Kϒ�3L��P��!(���P+�\����6+ϵG�ƪ��Ѧ��Q�or�������`��S�J�	A u�9#�5W��c�K��*�0���1G�U8l}̿׌R��L.�ھ�j�p�d�{���O�(���1)��k�ۙĠ̓�y�&��HIVj6\5N��'ol�X��P��3��F�3�V}W��czk��F�y3��c��;�cm��,2v\0����~��F�M�#�ː��x���H7�� /hSY�_��8ҥ'�r&)}իqb�6��Ц���h�f[h4W��&.DU=���s��;:_�õ[���+��5�B$9�×�D :u��
���n��w�ӡ�TJ1�OΠ, t+�����]�r�6��'r��2����?��W��lKQ_�l4��J��V�V9�Nq$�N�Z�=�f�p:�F�:6_ʇ�nb$�b��7K��y��Jc��+
��w�0]+qcD'��(��(p	Y�<Ρ_��7zM�%�4�0��+7��������#j���9���+��k)���Ȳ��=6�N&�	9|�O��9�>��eר��_v�w�{;X*=0��@�%���]���z���)�<���_t�Iu赑�VH���q�8]���ܕO��Q5d]��}�ť�[B{rj��7Ѓ��_h�j��y�Ƶ�߇J��*��~>�`wƬz�Hi����m����ȳ����{���]� �=�D0�f.��L��lV,��J	�fe@�6�m�4��<��z���~
[	 �]�j�)�|�B�	�����(��	��͟Ib�w��3�W3��I�[x��};6�u�,F(��d
���N�x�p���+!���
/�9>�ە�>Fe�o�<*Kֺ����]%�����m������-K@���ҁ�A��m�@�z��U6�zG��D�aw�r�.niǖFy�ir��C���fw�	6��������O0-`�" V���Y�랁R�V�3�R��Ŵj�ɔ�gvy9����P<43TZ,� ��Q�L�K�!w�EP^AI���P�u �=5l���Vl]�,�ɵ~<�_�	-�Y!R�°���k3���Ŭ�O�ʛ%a92𝅓w�Y���n}�ѻ��Xd�rB?P�{�z�F��$�4��c�K��k���^_0޾��<�"�whk��Wl�k�Ґv�<� ^��qU�<Y�����&�u����Rb�/~�T�i��z��������ˡy��E�r���y�7үy�|�\��
�P+mZ���ya�"���XL��@fC�Oi�c�ٜ��cn�i�bU���\A-��F*�/8�>bj�ІI���/�٤��O,�+?��Y���&&�+���m��ệ�5�PT>%q�*�c����e~<5�bw7c�A> V�x��vQ����ql���E�$�����^nT�EK�#C���m�Z߄e�Tp�;�׾�y�_�\Th���Y�u��s�2J�u$�:yw�ϕ��dyGtY�+J����N�� ��'R��k�"�ܙL��vn���M�B�&-�$<�������ů{.5\�H�N7L�5��^��(t�,Wb�D�nR��C5��������l��vKO�z+��fl��x���T#�QT�z�J?��1�8wN�e\���'k�]�;
�dK������_��̽�rKW&�],.ۊ0������� �jg�GH8K��\���/������AB�]�f��e�QG:7֏��UX�
Zw�s����	q����f�)Ui�T�F��d�;��鏏�Hy���+TU*���������`PF�s�0ٖ3dy��
�%�������"Nc4 Z��iZ�KK�jUӭ\dS�9�C�,���4�Y�=/tA�B��2JP�:��m7soTc�ߋP�~y�v���D�������=6� �[	�e���07� �D�[���8�L�����E�y�=\�Mٴ��9�6ȟ'3����P�ڸ�>����r�*)`P�dqf/*������d���~M�=���a�S�[Fa1�\S/��[��iC����X���k
�6!:��w��7N��r���#`7�L���ݪb2��Ѫ����]MpK�S���4om���%�3��"��Z*3����]�1~�+%|�A���G>�������Ό�d�z��
aN5������z{��JOS��#���}Mr�ο��(�'ȹ%�O%���P�1��]�������k���!p�:�����i�Z����f�:�-D�bD�!ci9[5�������=�Z�����P�xxڵ�%İ1���I� `��X3!�QZU������%�K5�<�����iرV|@ʌ�^��ƾ`dsx{�<f?*��qf�6_�{w�;��z��k�<CS�%$Ngv:?w�\<���G�<��%Ӿ�;C�N�X����l���:��CZF(��'���q;�t$�;Dp�����곣e��H��
�<�w�Kv��7�W�p��Nxa��mGv������SX�a+��I�5������K�?n����2�J� ,T��)������Ҍ%,�ܼl��A��;��n�4��~�	�]���� �Uc�Rpo������.�1ƛK<���7�D��w��&C��c����Z|�~h�v^C�|����M	f��N�{��v넾����!k��fO��o^<$T/%��Re�|�-*E�-�ۘ��Y	^�7��5������G_�N~�h�a���xn���zDy1�*Yk�Y�e��-��T���{�3G�%���~q���#u_yX-��)IP�Fg3٘�Sm��$�O����h�n @�21���"�`iy2	�~4	�^!��Ϥ/0�KQ;�I���~mU�v��Ŋ]���Ti�v~�z�RY��숲ENy�}�����<ֿ��]`�[��B�*2.w z�=x���AL%�A�j /R������(V#X.)q>�bLHp 5�+Y��>�W1#��w�^����8yD`1DC{��U�x�R-�ؓ�>R�����Lա��+�{�ݴ������MM�k{JI8��H��J�1&�'� �D,�>��P|�.�3����ڒU�h >��Cn
6�Bsa��/�ߓ7JYb-Z�_S78i%���I"�@V�΢z�sM�p��6�Ё���u~x�3�𑲣(D��,&���~52�\;(CS�uF�;V�6s���S���M�p�䛯V��3���O5Zb�����E��=W�h����	 ݀N�=[S����+�#��j�Q�^����:g�*Bz�����+)Mj����}ù� ����Q�;�
Tg�D\�7�B�c��B�?�U.����J�j�s$:L�ӘϴCS��<b�s�4�z#�&3�9=�F,���'��̕��d��ۦ8V�b
�	$�u+���	�9�ˌcŤ����.�5i��~p�Ǯz�?���926;rٞ���G���42K5�K�{ڎ{�S�i�*��FܚK 'pDS�3���c���3��!:���Ю����1[���b��5��.ѭ��3��[ӓ?�R��m^jh�zk�"7���[��:��L
Yt6��c�C�Pz
'���agn}��!��,����
i���7*m]`��v�������]bo����R�����8Æ������b��<��3�����W�6��淺�%륗2���|o�Gފ$�8Z��� ������l#�O�\@�	Gw�g�kb0}]=�'.������Ѻy<�U��؛A��\M'TߜRg{?{u1T|)�3�3Ip�!,TB.�Xm�d��q ��7&�'��8F���}5娯�$H dR��]7u"_Bω���9\8�� `RJwR��a��c,�l�s+BJ�ѵ\��}� ��3�!nz�&3���&�n��&Tʌ�i�|���f�d�����`�22d�|%7�Oj ;@�	�b(3X|Iو���hf)y���w8�$�[�~�Zp����Y�4��)c��p�d#���u�R,��r�9{	�mt���ߋۑ�:)�֑3�M�ˎ�7�H��yX�.�ȳ�2��
R@n����o�T��(�/��r�K�p�}0�?f���5r�n�����B����Rl@#%c�񌗪SKh�X��ܜi�d�:���%��?��
����>�|�.��$��h���{�8'~�3�]��5�Fj0��]�8�d���}H�ڞ�՝$�]V�I_S@�cpsS��������[�k�n������̗�15K��z����s�>�����l�v���m`�
�&<�2Q`�&��T�����0��_�L���a�*����؍�� zO�sC4"'�ֵ��zn~�M�]��W��Xb�b	ԧ~�s��!9�9r�-܊;��i�;�ꒄnU��
�����L&�͆TD�M{4J�[�$4=��d�t](P�]L[���� �I�����׷n�ђ
˹`�OϤ���ĥ..e�S�#����1�c�b��ぶwD�5�������UƉ�Ǯ�싁G�(�M[�-A���F���|�Z��d�4��Xq�(�
l{�T`�	���Ye� ���izN�(��u��U�%ұ�C9{l�4x1�նa7�b��N�2ƼE���_������`W9׀9�MT�����m���)���@�?��9��eMw��B3�y:�E*I���5�}�� ٭ҽ����[���>gv<�'��)��� b�|:��[��!��دA�������_���5���rc�d�Kz����g�n�Z>Q	���S�:<m,�Z	sJ��g��=d_a	�&۞Y*�W���\[�|��@��OC�zl����4�Z�!ص+��	D�X�����;2�6��*��O_�>0lL�[,+�)��ܟ6Ew�`<,,���}b9��B_W0mM3�3�τ/K�Gj��;�-1?h�	�S5�{�.�Ɨp4��f�~3��N�?v�S!k�ٮR����_��A�	\�qW��E{,-�~(@=�6��%(����{��	a���Yx�[5"��uO�G6�m1� ��fAO'Ʊv�� �$.�s�op��C��T�(7�	��vň}^ƴk��BR��V��>�R�㭀!o_����y �Wl^�2ͮ�1{�Y�5�J��%������V����� ���������Բ>����H1�rU����h�ژ��~1XG��6�$8dS�Vcg�I�A 3��	���z�x�JJ��e �Ü��S^��G��U�����a�*H0s�io�Rx�!e� >�p%n����d���$6��oN�w�f�>u� �����1Cֆ�ȋ���o/���z��N�������/(S�~#��g	0G�	��I�y�:v����ϘCh�
i,�$V����z}�����*a��z��Dx����;�.�"�FeQշ��@(:nr�-=;�Z�����<-qjikW�!ҢM[E�}8���ý����T��>���䠎�Gŏ��oP��S ܛ�"e�o����J���Z��%"�ܷO�O#�i�"�:��I�U�w�_���q~��b\@�i?i6I1�N�p^�(g`\�J��(^�ǩd��ISI���!$r���՟��W��e0K{��6F����5I+�����|�W�?�T��h�'���`��A��S��]ڔ��\����gR�hɛ��̰ @���A@v��2a?�{�2�O^���z.���Q�|%�����M�h�\*��7x��Ć��&Й�։���D#��S��<	��nЁ�_�v	8]����>�Ju�e�c���C�>Z�{ʛ_�����bđ	�a�n�<:4�|��i��U�z�g�dg(�
�����Dq��-�8�5
��S����^?��x/,x��N�d��zʴ�v�n��2���P�����[dC�����8�˻�)��ѿ��{�_��u����q�SrX1EP�z�|&��׊���� �p�i0�>:a�����0�0�E�\g+;ٔ�8f�`�.���,X>����{>����>�.�g��T]v��I�2̎��-�J�q�|{>��d���1=����1]7*�y
6+x%,��俺�>+ ����U��`��69��c�L�P�U�'��N�C��ZN+��G��<˥�݇����w�p�9-Ś�g��}7>{�.�>4�_�)��hW�4��xz{����im7�;�a&="9$����1(k��ڔ�Z�M>�YR�������}�`H����w��>>�X�6�/%��'ew�|�17w@�*���U2�	NdNm3(�Q����`@G�|d�����!�ge��J�p�N�>�O����X	}��l�՛�q�.�5"��}vT��R�OH�
��J;�b����m��~�x�R��{��|U3���*�j�y�< �$��X��W�&	��-�S*8��28��@*�@4�K&����Vh}O[��`����L�va�=�K��g.ED�B�,�1��i���m"?@Z�i}S��!`s�Y�yA�O�>�<��V��YY�h��w�e��0��z㫑K �lߩq�e�tm��=�9���+i�=Ax�\��
�U��AS����K0����q�7$L�r`Ǒ�JqkG��,�j������L;龠7��VD��q����)���Wj��r �s�=�Đ���ʈ�����l֎���&�>J]���n���8[�f��Nm��|�;^��s��;�Rm�@vߌ�2��2�ݥ1DV[�|U�7��]J_Y�����S��YN>c�.���#	 u*�[���vwb@�Es)#���4�X�l�0j���K�g�
�f��(��� �:X�HBuN��Bk�ɉ׬}˭w��E����b|����ag��&)
r�U�i�rH�M.�u����43�tKF��s�o@� �$2��x	_'���ś0R�O��@*;>�����0��;2�X<�9B�.l�\I�����Q;4���8�,Q���ǂ�vHDJ�&|Ґɼ���E�\��f��p��T���]��^#��=A�����K䌺�g��I��@x�����w��lA72��@�N��͔�0�)�s�g�hFy���1a��@���[��}	>�*���75�=q��Ӈx��k-��g�#:���$_����҄�xNX��ԍZ:��68�r�%������Jwd�Y���t:K�A$����9� �#u�pj�I��^��2kX.4|h*G*a/m�|?��N�l1#;���B��4(����x��� U��� �s�NнP�I��"O��E���]�8Z��q-~�m�R�=�(#�Q�!i����
�v���_8��A��	�JW	L����+:����<k���l�<X�a�"���FY9�k�`��f�m���Â�E5�ׄˊȆr���BW�\��N쉗� lk8�]
h��w����4�A�F����ck��q��`�e��WeQ��o�5��7�[ZZ��H�`t�d�WY�Į�e�G�^��Q��[�)��:�鸩u˿��J�U�3E�&?|��� �*z�v/d`W��k��#$��(�x��OR6�J;
T~�Bl'?'����S������rwFNoD5�������Q�4�~x���ˌ�����q�)}�!�̳��t�z��L1�.��V����2çB˗�K^��m�!��l����$�{�{]�fp�b�f�=y�� �&v�FyM(t��׾�!}w�9%��!d�yZ�0ϐ���?���,�@��-g�G���
y�`�K؟�A�v��7W-��5XB��s�
��s�3ꨈ��+k��H<��vu
]LvE �[G
�¶���|7�+���m*yĠ��u����+J!���׍��*���J�'-#	�&��4F�+�\�lcP�x�o��7�Jm'8
�ٚ��t��D�����_�e�~�����b�ۍ�F��#9�B�Qe6�ą��=R�k����7��� �:��GSR�6PO���%�?�6����$�E��W��*;�#�rN��wl5�s�{	�b����KF���%Y�&�A�`����T�m�
�执њ��)џ��j}8%T:�@�]� �;��KN��ًh$`�wa|��&�w������w�)�t
jw1��F	���~}bnD�SNl~�to 0ǳ��ͥPt��%��W
������B]m�\����-~-Cm����̈5V1��7{o'����S�Q�4Mk��j|���}���hqNg5�����FS��匴%�._�![��I4�d��e�gu8B8;
{��T�do�\C\�@T�zGЉ���0H��@����z�꠱Ј�h/:�!..��X�Cg��׷ī�N�6~՘5>��5rR��lYg��
#���Ǒ}���x+p�e�[�[�g�w[��H��4�}\��
vU�[�� �>���s��^�a�RR��J���f\�~��J��h�T
N�2({RJ��M�Jt=��/P��y;T"�>�q�?nRv�x�g�N'&������͊�0z��'�χ��v���`��n���yE��R����2�,��S����d���D;�m\o��_O9�?V�J!��3��]�A�3�H@�qhq1���A��*.���R@R�F�>�T�鐫3>�"�''Y��뷞�\ �9igde^�S�N��-�������y]��F���z����K�ZB)�'���6��P��aJ���_���m`r���K�+3.�4�������v(��F���Z� /�#(7���4�Ț�/I!����J%��-�� <���o@�2�E�s%��Ռ ��lD�r�ܝ�UʽU����\�p5r(�ߒ��i�[�Vy8��7�dyi�0S�Y����S��Q@�b�[*}��-�oko�j�x��:�_�b��	l:
�%��J�A%�n�jG�״��\N�5Z9]�->z��ï�Q��iL��H���/�*��t@�OA�+"��2�zZ���&2x��j�f����Z�y�A�˶�H��Ӏ�N����3���F{M���^��C�:gW�=_n�A��Ϛ)W*�����k���Es����*��ևN��.�25D�{7�&�@�!m�1���^����gj����w�+�ڭG��${d��*�#���t�0Nl�e[�
js2"�,��KnzL��"V� mx@f��\�V~5C+o鿌������u�q�\Ōeq��M2�s5��S���[�����~��5�RZ�9 X
p%���\?$���
�3m9���W��B��[(�H��e?�leˆ����t�j~H�
O�����8t�}�v\ �ݒw�k���2 9M|�z2�.}�jO(�N�����׻ׄ�v��`� ��bn쯢j����00c�K�u
�u �߮-��k�X��1S����W]o��/z�+�=�6����s��U;q��S�0����U3���#��bw&���=�%�+Ԥ��U;�4\�\����Aރ�R?�U�8�t����˱A��E�|Ҧ	��� 0�#V@P�x�=�mZMQ�b8ow�j/΋�zT�M��%�(��E��y�u4����P�n���в%[Wr�^����/��i ucm���ZO&y�"�Md>�Z�2��Y>�x �Z�3��d*�����N��ExW�2��Qϛ��������0���h��ׁ|�j����1��������^�s�|!�u_���U���{3Мv�8�XQ��+�;�����' ?Q8K��a��	M�5��6ד�im�\�p��'�B��&K��
�v]X$|�i��N�8��|�����j����u7`!a�#��Ɏ��ʽ�T!�`#.�C��B�z&<�+vS�|�4���&S����7TmǸ��!җ��KjH�4�E{Ǭ#G�R�>� x��!�A���5]T4��R4�%��+�۠���2 �vT���=���<�R��ƌ��Ѫu�B��hH@g��.�� �p�����Gٙq��^y $E�!٪�2�={�?c$�6Y���},m轵ǒ���E�S�X_�wl�!�Έ8EhMl��+,Vt����'v�7�B�`j⚒�S!��Y��uF�&ۜ����ޛ���l���kN^p^/�@7�����[��څ�c�*`/<� �e��!�X�D�)e[3k��׈�
��%��uB`Ⱥg=P�b�q���N�樫v��Կ���+	��0�3٤�4��k�����Of��1�$�����}�ũp�dr�_��b^fq�z}�Ụ�G՟�ճ�+�o�-{8>�Al�0�C>Sh�4��m�8+\5��/��x��~�J�w�d���4�F|�b��e�|�]�?μ�H�cX!�m��
BqZB��}yx��{Em_�m���2��:x$�I�s��r����Fe�E'¡Ѝ;3s���٬�� B{��B�ڶܽF����tG�O3���Eϡ��	�e�Gc�4 �F��9�&#�{w�e��qR��Ϋ���~-vxs�ڄ�^��5\�������4�t����"�~�oZ�DT�:	~�<g9A�M
�JM� bVz�	-#���X��#���tSs<��)�ns<�*��)����7�'$��x:�I�x�l����-@d�kz�L�w�d��&:* ��J���f�BEN-u�TC�����c�20C��HԫU����;�����1+ H�y�l\����|sZ
^�������t���f͙WOM�r�#�@�)�x�ޢ}��Ѕ��iB���x
QCc�͆?�X���?Q���
����9e���^g��dZ����%��!��)���r�0L,�
#��bC݌W�.^�'8����NHx�G��6_6 ���s(q�����H��B��0/�K-U��"�����>"}��2��ÜF�pY#Z��� '	��Q����>I墇k?�p�VH&sL{��T�K���מV�UVo��dZ�~��@����^"bT����֯G4�!'�3����&h>)��>��s]�ύ�~��Xi�����Q�M�j8�O�����8����� �:����a��L�)�7�ݵ�ptt�E��)�@����Ǘ?	tL��"c��[��$eXR�U'zL�`�}X�2�1F���7�fqLp�(�å�u֙��׋��	�/� ��bx|�I�A�b�=�oT�(}��|���[H�RG��!+D��9�r�e���mp�����7�z�;K�����V�˅�B�0�3�PO|�ZK��ơπ�pIƍ?t��X����eqU�ㆹ��S��<A{:�]ǳ��|����k%&+RKbģ����K ���Ђr2ܡ�T5�_��z�&ߝ?��HH��k���qb^ӣ�N�*���D�����-�a�ΛNQ��1������"�H�hhE�<��_�*���a�mv�L|?�'�p�B�C=�p{�t|S�^U��9�`�
� G�հ�T(u?��" ��fֆi��~��w=�.E�ԏG, �忀�N��gl�>�;>�m5x��~�Q�"�@��#[ܩv��������s��*�Y�^�����ּ�� ���79�BB3��C7咮�%x�$�RJ�J�Ih���J�V�r*�Bk��Kd|��"Ya0xo�㘎�)�.KM�s�� �m0tS�юM!./�Kg�xc�|3[VXu�Ѷ�f"vK�E��[Pj�Ffo�E�ip8�z/I��X:�iͶ��Ƽ=S�k�)f�`�$	�[�4G,�ȶ��w��Z�d,�K
���{c�*Ӹ���y�!�Eb+��h��B!��S�o�	���wua.�`х�[�b�>|?������|�|r��Kzp�:%/�ྗ��[I�fu<�f}۞7w�0���z�O\��=d���y�0��-���X�đ,;�z�g5Β���ᎾG<�W��t������&=z�X"YTB�����"�x�B6V[r�������b]�7n�-�z�߭�ӕ#�6�l:��X��B��i�7���w��p�j��7�U���[��;�	��<ֽ��a�]
�=)؏�[[(Zt 4v�)iȟ7��Ύ�S\��@KB�2����ğ\;�8��'L�D��Z��\�B��))���8�=��n�0I�)�V��V�Nwf�d��ݰf��nˡ8�\a�	}Ļ~Jۋ�����N[w�BB�G"���������p̰�C۶��aMCRnl��0��t�H+�6����֮��2DyAnF��[g�Ѓ�"���z[GX
U��F�"���N0�vB��=���P𪇩	�G@�Sy�o��n[b6ծ��"�1&��f�!��T�˹�QQ�a"�3{ؗh_T��a��$���J�F�	3�H������rw������ؓh�U65��<��� �ur����
�xx��\1	kǿER�Ԋ�A93��.3�f����V����#��i��y�{ip�ј �/�1�C�/KR��P��]�)7��6D�j
�]½?_0<\���a����%���#!�е�3g��
l*�}q3��"���Z~�����.9�����%:JQ�~�0}su^�Vj�W	!����I��ye�&B�W�����q+�JV	�
�Y
�A�O�I�*�l7��AZ
��^�,�V*ű����M�)�R���Q����; {�J����5��!#CNЃF6�V�	�iޒP���y!��u~l��|��aV�֒��$�{�"`#M�5�����FX(j�e�;��4}Q�\��V^��T��o�K���{��	����P�k{G�n��f�TU���ㅠ4k� �I#(d�{`&�=P�kٙBut�#91�s}KAH�I�";w2�����\}:�	�k��-�D�:��ֆ��hi8lÊw�J�����)��	�݆���@;̂GoF�ɂ^��/q�6e�q>C̳͓��ͭ	Ӄ=�G���Da�\��ń�V#��Z�~���<�"�{5f��)Fz(�L���ھ��P��_x���[�w��D|IPj��1��lE7����z��?��:��?�ui��2�N�V�cT���jpBr3�%�ۻ��y��)���aO-��&�����g� �q��r�2�dٮ!<�Bܝu	��B�Pm��F[��#,*�/��wKhP���t$�E�޵�vW�<����C����i��TrQ,Ɗ������'q����i�4%DA}hϨW��|���m����>�;��pC&��i�a���. 1�P�Q�C�-O��A;i�IG����LB9Q�ְ�����Ȑ[
H�)܆_�_���H6��DKy�)_�/x��V� X�-�/�����;��Ty_����N��� �s˩��0��hhn[�y6G*�q��Mp�$#H�po�+�r+��l�o��J_b�P2�Ծ�g2���K�>�F����ɜ��[�7��h���q�9�)�|�w��)ˠ�V=a�����_s�����������v�e��R To�˫{�u
�Ew�o����j��>lAڔW'�e������.�ݴ���q��z��}��[�ԈO����T�ܑ�/����8Z���%s5��i��d��H��U[��Ĺt��=��y���)j��p����L���0yG�i;o�t]?n��xsrmr��+W�f��Be�S%����iV���>��g��(��&߅a�.D�kM�:�5=����z�<�����4�*:Ǽ$x)o��`�D��Z�����d��1�^�5�^�9g�'�P1]/y��a�`�[ZŮ���6_$T��)5V�.�V�5���Rz����-{�v���0Bw��T(�Q�*����&�RWRcd�=�V?<��	��;VTO$�����[�-�j	����M1��m�������3��E���Bӻh7��c�&c��`͜��F�Ik��� ���V�j��Nd��,%7{ST��̏P�"㸂m�|���(��{�"#���
��3-Hh������<�U;���ޛ��Q�8*�P��M}Z�Lw=_zv�P���T[:���]|�Bou=�֏��b��;�I��5�XRG*��i�����7�M�eP_7��{�JTα��/H�l�#��&�&�V�=z I�}��^����@������J�4�'�BX\��@1�CO%F���}����d�M�_7���kB��.�s��"�盗T��l��ԩ�M̈Es';�4�S1
:��N<�Z\C�8R���$V*�1d�� ��5��;���Ky����ө���Pf��=n���KQ����b��&�mM�4�$)�2A�����b�d�\�j���P�����ZF:=oG#��\��(��#�|pg.��R4���>��`s���{��&��D�����V⚟m�^U�z��3tV:���̧���J�}l~���c��3��lQ��_��2
�^�����I�Mb1�A^����/�\nk��8L(��%v��(H>(_�\��Kَ�Ӵy��]�7�iϣ�)W�����w�;gn�_��"��F�#��28���qM��-�Sǀh�&y��AMv&��^8,���,���X
�m��[���o,�!�^��۫�Į>gc%����7���eUm�E����8H��eaL�\l�Ba���7�A�S
������L�p+��dzZh��J�2�I����861H�V�(ڮ��i�ʓ����)=�9����8����/1��(��fR<c�F�s�5��]PAA3��I=��c"m�\����61��KQ�1R�ءP��
��Ɇ_u�:��hu	��O�,�~�g	ӑ�O�;�|/.@xn��������$��1�E��E�}^Hͼɜ���$vw�ڂW*���p���B�qh��13s�4���(G
����]�v����[�B�*㼚�@D�������+��T��H!*R� J�Q8�&ۘ��y���%X�1�/�o��a$S1��tkt¿�e��;Cg��������l�,)V����kL_g��d�V����,?���iE�ĭI@��W��tɍ�i������n����o8��a:M�(�b�ĵ�(���#��Y2=��@͔6��ڎP Fng����w��g^8N\�W�jSR���?`������E d�侽B)�{C�8���i��U{��y�z�˿S�y#儓��8��;�@Ȁ���gH]�x��[�%�]K��^&h/�����+��;��U�;�uk۹T����B/:/O�a��7}Ƀ>m�D���O��`AB�����cǙւ=h �Y�
P���r�k���u��#&��;C��3��ڤj2�q,F_ޭ�=Q-N�*�����n�7q�P����#y��NE._�s^D"�
�z� ��b���g�U�Yk���ͼ nY�Hʔ,�v��0;���;+B`!����!^��*��j���0�d���������v��\S�4^�/��]8�t8��#}ٞ@�N����+"B��F��'����E?77Pɱ��() ���h)Ï4��/���N��E�O����o�Rrb
���b=�D-)����k��Hy=�b�B3�%D���$j��
�7f
!϶�&��|4i5�����9��7�[+0����Y�X�X�{ �\��$��aVeݱ=�P����̍���||���Т�ǰθ?��ٳ~�G���S�+�=?�}x�R�@8Xb��v!���c�}P@jN��J�%}ۜ�
7~ވDL>�Ģ�GJ�rV�Jd�������Y�LAb�e��p�e+� �I���O9#��Փ���3b��0���ǸR�_1])Ԙ�{Tp�F=���r�b+�rN�ٴV�HU�}:�Â�3��Q�e}ٶ�ȸ!4�,[�ru<�oa���/���ӫC������fA�_��lF�[�ِ�B����	-��P����SO1� U2��,<��Sӧ��q�3�PX{{4?�&��qJ�}&��Qx9g
�����[�5�{�w�N�n%O����t�(�E���z���X��G,�X�숬�m�����L���l�0��|�)l�D�?�e�}7�A�旛K�z5��|^F�⺓a�����?ʥ+�xj������
�ӌ�Ԅ҆z���p�#tV8��rO��`_��Xa�ll����U{�,�.B�A\�3iv���%�u`C�*����T��ϱ&�d��yYn���!���آ	U�<�潏o�?!?6̼?�ǘ*�װϬò4��}�y����t� /�Z{�,�ed>��c���t�ll����^E�:\��Ӗ�^4�G��f;�z:�ͪ,�~��_�������J�#G�#�,���<D"�⯁�Ҳ�Eyˣ��@�K�n�|'k�\��q��++~F�w�s�F�Y��"c���^�ù�Ag#���o�7��s�K���!��{��ઝ5:�x�C�]\0��}�I *�0�f���~1��Q�g�ϒs���=��*�;�R�İ2ɬ��$�	q0�(��I�_/&��c�n�q��%���[�y���V[ɦ�� �;A��ϟ'��^��cg�7䷒]��q/��r�u�)$?�H� �j�]��y򞂧��վ��A_��&���Ee?M�����g���E��c���UwA�x5��MV[��GS��=���ھ<4h��l�%�.��4�����9F�x�1�g�Dm+Ǳ���1��w�DۮVY3ٚ��i��K���j�A�\
T� c���$~/B���#�<�tez��B��r���'w�{�5���=&���R�<��t�~�?-��Y�1H5���-�79��j�RX(����=�#G�{�伄�q ��'�x7CH���Ê�[4	P��-���!�}����%�)RX�]xt�!���5ȉ�tp՜ى5�@,gm�͏�u5�d���]�((:߭ė��6Uw��~8���i˱ǆу�M�	Q���
rSg���	gu�4��˛e�I؞'��­1F#Ҵ$��jS�M5��X�f�[E��v`�M�=�*�'u��8s��m�1���ŝ�+j�ޱIo�e�˕4a���/"a�_�����D��5�Oe�3~5aT޷��ȋ�wY__�;<��r�WJUv��C�1؆�_�M�_?|��ː�4LɃ�u��G��E��B�6�F�s�b��'}s�{�o�a�f�6�-Ǒ��M��/�a��z�5ʄ9�R�j�]�ْ1Ä�6@�C�J.`�x�_!�\�t �)��k@� b��A��<�s�h��ܢ�P��	�wg���L1p	�K�or�R8�P��CUL~�3���a�4o��x�"B������L�6�pt"��ׂ�#��O�4&UIr�>J͏��j~M9�h)0��Χ��(�o�k�+.ȬT��˳d�W��Yci���=��/��?^�C�:�	^�R2�B�E̬���(��}��Y]�y�Ew������H"w�d�y��k]�S�*裆�֐��Uё�Q$�3�dq!D�R�>�;gb�����!��8<�8l,{qZ�1GB(�^���X���U���A��~�Cx�D��"��8]3�y���yF�3��^�@��F �R�F�r��+J�(�A8��w"6k�FdPB"Ⱥ�f�&��*5⻓hf���s�9g1>0*�	mB���w�hRNv���j�� ���9ͷqǁ��ߑ]EPoi7';O�o�f��_+�&t��Rpx��}����N<�`�-^��T�A!��'Z��XI��̽^#���X�$ڧ�7ɢtēE�Pۡke�j=5�S�T&��a�dp��@�O$}��Nҷ}�Q�rO#��r�띩p�ݗ����n���i͏+�W\�$��+x��D-���O)�"��:��WU:��xI��c�#�'��
������J������^��9���[�_cHʧ�,�7R�_�� Dbé����)��hx�ߍ(�u4
�8lJ��*2��llx��r�`�3�0w:b3���C4�襌5��`h�Ar���X�*����)����\�w}��G�Eױ��͟
�"��8P.�����V*r����� �B�W^���〜`D󋇄:�1; 3�`����>��i6�m:�tx�0�2_�����������U:�@�"�f���
W8QZs�x;p5k��ճ3P�0�$�� ����e�/'���m��1�;`�J�h�w/�E�]�TԆ�`]�X����>�E�K�!�蹕���x9�@7�:��l4D
����d7:���$�������qA�evwTH�D�}J0'݂�Z����'�硎�+<�=oѹ�i�o~agP����u�N�%gc;��>���û6�D�$���
J���"�D<�>s���I&�o�%>�Z���Q|8Y~��r�RM$;*!��h��U�L�!n�#KT$�w]���a	�,��B� :#_,Ag�*���'i���/ۭ���l<c����Կ,�,*Q�ƾ����ɤ��	y��C"��`���C0�7��O�d��p�q��^��3ƞ��_ ?E�u��``C�lucpk�I��n�q�"�/~5�0[^ک�ǰ�c���P2O��i�B�N9�6��I�4-�a��!�}}��B�E�iS<$pm%"�<r*�6JP�t!��y3�k�_+tj7��g���5!���:�O�x&� *���Y9�wK���E���AvW�i���c� E2����+�7`]xݾ�U�l�O�WP;������O
��&���X��^+OW���,��.6=���f9"<�K����j:����?Z��_�����Cx���������%53d�e`��Q��>\hW ^ߐ���.�b���I��%��!�؁GM�`<T�9#b Bs�E�T���8���(Z��B5�������/�oU(2�;�U8�'��f����$ظ�6��4l����1���E�N��&�����n־�"��*�)���M�s��).�is�N�*��~�ɷ#k�4���ovzE-Y��J�j�h�򴘋Ɍ��:+T�RIZ��G�A�%_A(�����oB6�����D���Vg�����+
�la�$j�J� 7P�w��G�c�?���I�����k��W�����+�k���@�^�:���e�҃�[u���9N�� b\�2*�rZɂj��W�\��c#��uDɍ]�h��Q���)�"v���kHN�:T�|zՁpH��|b{��c@��3U#�Z�!�X�R�x��p˧�<�j��o�p/8yp��K��캅�ly�����Q�
!xm���zRxbS�\��w�'����4��P��P{��[94�|���MO:㱏��hR�$��?���q�ې_��`��O�o稏1S�S�X�:4��U�b�e��0{s�N��$r��h5 ��{��PT&��)��#C��Eͨ�7ک�년�?�R!	H�?Ef�f�����V���3��A/O��"*Ч!B��U�C�J�9�x�B�;��p�Vu�@���[)�UV̉�<�牊��$6�H��Z�ab��P"9!��� -1��G:�ǹ�z�=���3[��^�h�<�5��޲�^'�'���Ӿ��*����2�.���~�����uJ�����Qx�B��������k�&�cۭ���IC^q{b����x��4o�g(�̑�Ͽ�d7]����΄`c�
l��A_�5�B���L(7��o2���-J�-ev�6�)���_�ƙ:{ igZJ�UCE㭦��V���:K"ʙ:�}���N°�۔uq�����w������a� �\�5	���N���ɢm�������'�:
�#6tpI&����(c���ǿ;$�̬�dh�J�l�q]��T��cἍ
j1-�����yS��%c�,c=#����Id��F�F��q,��Z��{ã�r��6�g�D���>��}����'��l)W��qp[u�cV�j�=�I��{�YM�{+ŋ�q��ߴ���Yi索2g{t��傾���� �W���IA����Q������A^R�2���ͦk��A�q���|��|e-\�Y�@�����o7�O��ҫ�Z˼|xޒ,�b�̹��oh�.۳G�2�u��B
S����>[�r�<ϩ낋��6�Hdу*�C/2؍�cS]j��~�*S����l,�q�D'2{���A��Ӂ\�@�5C�L��p�C�?�W*\|Be�5-��jx����`�C0�$�J4����@�Ϲd�L���ښ��ӷQ�l�@ݴ�ׇ�W��B]�'rI7��5�Z9!�:s����,$��O�~z��Յ����T�h �������9���Q@�#�E��F�i�E���PW��W�������������Պ`v�R�R*��$z�__��>AU,F�15:� �4V�>�	L�$��P;�x����'��(x���k�W6����3�ֱ��W���nkeh4��7?�j�v.�~���ok��Zm�� �"���+�l����xꓯh)˙g�(�ڟ#��2��F�P�* ��
M���-��
>��ө�r��A����l��e���u�]H5C��ԋ�X[��fF�W��T����F�DH�����J$U[b�ol%�۞f���G���n˻}�/�NH��)J��Ncþ&�֒�|��h����(q�7U9�ƖD��mmZ^�����8�[G�|хf	���l����B
� ��<�$�5
?���'=f�qA�c��{�ý�~���lS$�c4j�{���57=��['���oB�������ަ�צY���=��Ƹ�&+����z�.LnMo�0��-�vw_�o#JG��:�^ՐƢ1��Βt�P�J��=
Ȏ�\5��HzUA��
�`I5�h�a�Ǵ~��r�dSJnƷ��w�� ��ۗA�?�n�?s$%����l����������G�0�������[��F��6Bx�~S�O����u�ǪT��I�o>�C;x,�o]룗�e�e������q�N����G�����ל��5lm��:����Dwd�ܬ�S:��ȧ|�S�K��y	�%�	Ц�ϛT���X3�9�;�0U�`����2��1���&��3��ϕ��Fg\՚m�"B�b�~[ޕ��ʁ�(J�nD�������u�����O����C�H
6e���Q��.��W��U�H���='x��J�$И�,$ym!��ꃗƬDX�U;3\�2(A*x�ƛ��'/l.�T�U(}���5	�()j�7 B���a�}���;:��J# >�������TD	��.�+e��(��O�~pZJd.s�v��`!�q	�j��]�5� �l�N���� x[�q�n(>%�{Fg ����J��F�&��>ʔ=��Rl�u��'c<�	�!��k�!�ZCo�ST ��'1��	1�����������>P:P�j�V,w�-,	�Y<��Q�.���2�p�_zFfˋ����f_�:O���iH�-et5s]���e��bO����)��b5NXŰ�7��
GB*J�vJ�Ƀ�{�M�YI��s�hz����N�W�X��f!M?���7�/*���ws=��7H��qU����A�w(�P�f_�4۷���Kؔ��l�nlz��2�k>�|
�{��}���M�v|��İ��?8�H�FY�f4��C���v���G4����-���w�]���$��#�j�����s�h +� �z�w�g������X��T�kW�]%�,�e�M`Ϊp`��y����&�����,�Fݺ,?�m$���aK�ʝ�	��aHe�)bL}f_����cp��.D����|��l�`"l����$h�F���SD+fY�KC����!��r���)���ʽ�e���MK�{Z���/�%T��(���ÿ�nn#anZ�y��^���l��I!Ǿ��vG�R
�~�L@K�6c���n���k���� `�A����H(����1���u1��r%�V�tS��;EP�1�5Pa4�@������%�H���1Zr�4�A�ݛ<�OOܼV�~"(P�#3��W2aBf*2�SV�1H0�Kx�tAS��[A߁1��u �0�rH{�����x�G�rka�g	F�g|(�ٕ1]+�o�:��b��f���ߩerSĜ_v�J{���IP��s��	����`^+9+!;�܀�j9o�"�_T�
�p7n�7c{��^puƈ�=���5ħO'�C���6��.M>:J$�zV1`���ExJA�g�,$�.��&rr�%�%��S[\E��wX2��t�:,y���}�}db^��[���%���wG���Ic��h�~����Pc(�B>f�#;�q�ĵ����%�_��Oۊ���H9�z�����bM|	9��Ŝ*�Q����o|�0tI��*yKE3.���iE��h�;���VPh���|]�U�%��8%�~�L6�N�өk�����S/�Q�
����r�ai���jH� l�Mqh���l��&t��s����bv�]� �^��ޥM"���� �Hl�R@¢�O0�OkXo}���:�ݩ���ۈc�[T\�C-�ʧCd붨f���*R�Sp���G�"�; |�B��&���SU �.g�l�N��|8u' ��
�Zx}����z^�a��G+��!����*c�F*��	�xK���ۆ��@:8��R�?��o$�_䀡�v�u+���o�vl��8����X��p��fG~&��?,�8�^l����T4����ͬ?��(Hh��n�e�D�J��Ҥ@|�����D1�Ȃړ�P�:Zm�q�D��}�J	�R�}�������-]Z�J%�
�pM�����3fm�¹�w�����C'�.�b�J�t2Vn��Z����6���-+X3��S�ì�9�1q~�S<�͒��G+���h���e�ѽ��e�}e0�)&�`��O#�5�+��|�����a���#xY�	,n��.b� V���J�9��������T��R�K��g<�T���n�<``�S�gsN�{*yf|��a�I���f+Jkx��#t�t��T�ဍ��@��*T��1���.��(���5(>� ����$İ)3�O�;e�\�nn�)xz5�Ғii]��>NC�[��v�ߌ��.��j�]�;���υNȈY"�����#,L�2GU�a�tx�K�\jm���8�߱��j�k�v߶��cL�z��	�b�/K��d��Tn��m��/����m���̞�ܲ%���b����R��@뇹͆57���U������y3��j�y�����Z0����K����H^ds�{�1��U��X.D~�8�/)V��J'm�N�^��W�Q�[��_�o@�bN��ّ���1V�v��٬P�ړq��;<��6�	�J���8�fʩL�w�s�'���˽*g׻�s &���[��xb	%3]y������py�:���V��L*�~�����D�)6F� �+��ɭՠ,�5�;aP`H��v������N��8�6�yُ6u�/��l�'�l7ѓ&P���
���0�����v e�6JaE�`���ur�����w�mu�a9ir \�W�����[7|Al)����ҁ������eke�H�){�|���Kʗ�A������ ���Jͳޯ��H�~<	�p7��=k�.�?i�����L���������᠊�a�G$/R9�%.�D�B����A�/�I��;��'��j�)�3���̹�6޲�\Y~�h�mD��Ղ�#�Wܶ�AS��R�*��>���{i݈:ו�}1-�MU,�SS�b��]��Xlf�t�5m�d l�+-�l��'���{ҹ�R��FkL�Bu_ߠ`/��]�*!F�,�H�<��_�NO?�Z�n�>j
O1|?9l�ʋ�Ź�)��/R���`���H�),LEʵ +�{+
��b��_"��*�*dD���7A��|���zS+ ��w��G�t�Kw#p3����S��m���:��KY���f*F̙*�j����c��	��	5�Rn�p��e���u���N+>qHD��P񬿊 �yu��}&�����v�	^'��@��O�khz���>r�i�y�̫�Y���I<�n�|;䟧,���^�?�Y��	����6�=`���rkb`?[�&�芲]�< ���Q��N!�s���1�QB
�G������f���22j���E��dvF�f;��U�˒ɠ�9y"	 �(���ʄR�R<{(��Ǉ�&�j���p���
f%K9k�Z9����U4������ó�Ə/���j]�"��؊��u���<�;�s�x���~v2`	�Rm78���]v����������EΜ3Tn��	e��Ɍ0��6����Z��ȯ�s��!�c�ւ���>�57�����6�e�71.D��%S��cn"�n'��[�avj:쯀�M�ţN��r����;P�et��1iSn�~F�p��� �����qv�j��������Y�h3��Y-TE�8lqE�$�P�r�ϼ����Y:²��Vb-�,�9��f*���
H�g�z	�a��*�bZѐ{�D�e���L���I}������=MݰߡtJ}�������${�q^n�YD�L�])����"��0�d�_�Kk��	�lAՁ��䣑��r�F��A(�h����Y ��� �����D��Z�m����eiW��Y1=���1!�*��
�HC�:>D��qP��|���i�l ��'k �A�4���yz1_P9�-�Ǯ�G��M8�\ a�C��yq�A:`�H���C{t^��o/,`���^�t��#b���a4��
�0�D�2�7�)�:����1!�:�'�x�W�I?��S6&�ߪ}#Ϲ`�֣�5��pʯ �������1*��I4�������u鲘��1ۍMyI�.]��M���B�v�&�G@�䋶�豭�c��ϔw��Y!��L��4��:��Q�V�V��t/��5k��`+}BM*&&���I"�F\��mG8m��U�u�h��~�}�&�x��ǆ�aP���'7̃:N��vQ)a/���C��v {s����b�+Y��|Ъ�����)q�"��ECI��yc��Y�<= ��r#
S����`���R��"ٟ�F���P��8�u�`�c1C�^�LF�pF-����{?�h���8@B8J�"*�A�՞�X������ג�U%G�/m{�0f�KL�w�ˠ:)���Ĥ݅
�ғ�I(��E�����N.���ƐO�t`@���[��AԤ ,J��s�zRh�\FY`���}?�]/tW�x��w����&��^[6�!|��V�J�xŧ��)����\��Q��ػ�'<�%�r��~!i�������OB���T��W�}�T�l.��!F�3�*С�j����X���>�r���ɒ�!�����[��#we%����=v�*���vRf��	�=��7pP�֏.��t*�tE�:�c�;2Z�!^�Bô����gVSśQ�{���{�Y$�����w��c6��R��R6"�
�3��`d�YG��ae�`�@���1��O`Ue}�v�� �5��"�Ɏ�����4 ��/AT�Ȅ��hcB�����}
�D�z��(�0��Z-qv4�+���ۇ��;M$��?�ܼm�Ĝ�-Nުn����2�m���ly������d{uH���)�\���������1����V�j��M"���,�PM6�9��(��μs1��1���|�F�M�. q��h�d%��;�H\�04��:D :j0$+p+<p�Tx��mݫ�)�d���%h��X�X�'םP��;�LZz�G.��`'EZ��n��� ��r����!��4���S�
�{<��z"X�Q��]s:��;�������2����G�W�1P*�Z%�#�I��b�8�sR�JK6��⠎��&3�bO��[�\�?O+E:�x�J�1���IZ�(� ����=��������Wh��=���Ŋ~+��f��G�W���B��(���u����I��H�ߴu���ǄuZ��<�0Q�Ά���Z	,}��XK�Ö��u4��uRVa���jw'�O@{Ծ&P���(3����b0��S�
�
� �11U/Z�RCw��N�S ՗��
��y�e7]hV�����-��Y��	�X��N���v}pEA�*���P��8j�4�-�i>
�&e����3~Tp?sJL��*K�F�ܭ��V^$q��&/ �E3�ȜS�� �c�q`q�n��5��|����X�_�l^b���Fo�FgƖ���fV5�Ea�J��c<�KD���g�OdV�R�{��F��؜\,�M��kq`�f6]�`��Ш��6��<{�*������XU?B�~'RAh 5�����AZ
�cs�¯�(j^|DjNLՁlgX��M%1�z�?�W�m�w	n[�Q8���t֫�>�RO��e�𤢢y$�KX���^l�Ĕ��d�=�� �5V%���Gi�%^��c�u��ο���̈�{�.4�6��3{1:��?Ht 4�X����n�D2	�5:���R��|G�^��;"��Q�2�O��%B��1�㣦
�9�Ӏ���`9�'��"�yÿ�CO�(?:�>�Cs`J�:��y����UA��������@![�"�+��[߫g��<����fp���%c\b|���
��D ̙YO%�*�O|���e`=����N�8�{yָ��V���^k� 	7����>!��S^28�U��wU"��pռ�v!4��'!��A2�{+���*(2YD��׸�_N�ߟ��������NX�\���l0��$�GѠ������fZ���`����gW�~J�H�ןu�^R�P��(��k5W*�h�6*�!Ƣy�l�Nx�N&}�ZA�6pd�d��.H�p&������~�mY�E�h�DL	��@9-�3aK�0`���x���.�5���K�ס�6=�5����,Z�jq�s��� �n�/��$煜�ރ_c	Mŝ�&�v�Ĥ#S��Eψ��D�|�q�gߢ�-r7�O��f�_��|�7�Վ�47t�ͅ����G����vS�$Z��'0;3�9%8��e�k�"�U �nUx:L+�.g�$OիKa;�V���3��2�[�U����ѫ�dc!��G�1�,�Y��4�e,VڝSW���Y���e"�G�RJ	��f������mm�~jrt���4�'H�]�E�s_��C�u �E���t'x̛�'��n��g
�%Q8 m��j��������/Q�8=u�l;K��q�W�2�q7��b��O���[8k5��uQ�V�C($�fK@U)���au&���3Ֆ������=�Ԃ�dJ���p(������FΥY��"ڼ�%`�{!�V���|��,��\����t�&�����[��/N�|)Z~\���x$�������_�(�Q<��^�2bJ^i�QuQ(��f���2�&�Vr=<
��'7����*�6�4��vs6R���g���J=i}��rngϣT��1�d�FP޳ƥK� ��������@q�����\}x+�R?�p,�N)�ht�i�<�)�4�*��)�vM?��by��F�������F�˵քol0���8�s��.5�}8W��i�p��85��oy�J��y�dT��֥��˕��G�P��<KA@A��
ٗDi�q�*���(�������#�=�>ݤ���x�D��o��� X���Z�J�y7��G�G`G��.]�T�E8|H��S�S�S���9|D�|��YK_V��h��fRCJ
�<���A���#tr�n;'���{�$���U�R�\M�,���&�!Y�d@���X�f8%ӈF��6@`�f����ȍ����6�|��C��N��g�ۖI����y�eU �S�:�̽D�+0/����p7P7
V|].�qi�v�uaC�f�h���)��>W�eVf	������3���x]'&��R������������&�&�P�p��9�h#�.���䄨�Jq�z���ɘִ���@&�]�/�w���@�R�˫�p�ps�E!|�Q�S�0��y�|�F�f�j,ޜ.'�3[2��$��Ғ&\���A^�\�J��(���O��å� \F`��s!p�����T�%��E���Wٯ��레8�%m��U�M� �*��UǍ��3��x�h�D&��������J�^���$��}�[���@�e��X�;Pz+rXj�U`ir��2����K`U[-���b���Mw=;;7���{�� �����װ�~.���7���.���"�Su	Osh_�_�|���$���<[vk+����[a*��U@L��;'�>=T_���"R<�!&]nÁ��UB�p�=���j�U �=�4���M�i���BP��hJ5�(��}+�F�����qX_c��t�L����U�PW������D�&@L���N�m#t����A,G��yLb�"��a�FW�i7ۆ�xQɞ+�Z���Kۍ�u�T�|�Q_�=YP���f�~�>�����%y2�
�_�&�f�����qt�A�z�9�R��""6Mm-Qs�N��G�Z?ֱ/�,�v�͍��l��C%�
�3���P�f?8fF}Q�_�Tt=#��gu��*/�.�-dW�H������A��a�6F�D�=�Q��q�
T�Ctd��j�h�E �Ma$Oԍ��#�Q��KJ=��*�T$j*�rĚ(X���(̟���x/ŵ��6�ƀg��ن�[�\ ��u�tG �pnU
U�S��x�{O�82@1�I`�{�]F��2,�!*no;�ϡ�����׳F�#�D[q�O�n�V)'/ɡ�:J`��P��
��Iy|og"��_��ڙw��:��l5I��.�юy�*�Uѻ��d�_BȘר�s�	� �uyT�^r�aݿL���#m�����4��	��x�U,z�9D�h�%�]w��T����HP+DF��
���X��W�}��\v��݅(�g�pM��/A��\,S�y�XĵQS�=΢���%},L��&�����r��KG��N�Jr~;cω��K�X��=3�<��X�H��ol��������?��m#��$�!�l i�>�Ū]ꂭ)-����y�6c4�ݓ�t��ޟg���} J|nD�ѤN��D0w��f�(�U,����p�*�w�a��P����|��7����wP:�U��b�}�jz��p�����<�e�_��/>B�i%5�TK56z+Y)�1�Œ�� �|�){�A�w�$*Bd�\�����IƲ23G�ҥ^bl�F��~��Rq���P���8߅��J���YDL2M0���FaZ���Ő���y��y_�#��ί�xA�	L��uٜ_���D���ڕ�h��p�� QW�t�b��D�/[���H�,D :���L�E1�.)��S�-�4�Y�.xъ�	���f�@<��1��A�^���O2 �N��q@-�ւ)�L�Zw��IZ�ُ־ǣ�n�K����rz�;���+W�Qw�26[��q�/��
4b1�r�5Q��}lLa���*�����w���v*Ñ�6���EB����f�M��3�h��L�v��}A�C�HT�up��"TU��奫1s�:�Aԣ�5��C�o�:���
&򉸨g(�~;ڊb����u�Z�$H��yp����y�[/�*-0V���+3/�u�n��ʹ��`������
��~_�I}�bND����i�$Ua��u}w7�I��swcO�1L��8J�����B��@��:����P.k-�N����H��c�GJ�JHH%���s���G\���l*-[gH�j�N�Fr�6��)�@��
��P����:���X�hY^..��c�N*5��������dL;�K�$�Ia��%N�Q�	?Ȥ0#ߓ�����ԽˏUOr1���j����Xl����R-D�$ryG/�.�@��ª�ʔ����b�m���8�l'm�CE���
�I<�A��sb�u��Wԛ��ę��Y�ۊv }���:+�/ ��?�N�豕U��������ܰ0B�G%^ɢQ�-�hc�fP�]��1��B������{�.��^�2Į��r�1�l�0���K��D�� )��.����C6XwZ�f����9�E��5���6�/�������s��Ucۮs�9��q\����6�p"�ew�9+�5���m������)�f���$"K�8o�%��,�3Ư��?Z[�T��,t]��[�C���\7�0��֓{-85X�*{��6j	�G��*�n����һ�Y�{���E|77S�&B��(>�
�.;�YA��f,:�D�j����L6��.���ڿ�-Ŀ���-c��3�T0pڨ�:�^��1L�zm 7����>&{݁��C�|d���S>4��>R6{���LNܼ�ڢM�.�J���&�;2ma=q�-��=�����
�%I.�@�_xR_q�6H�c<o��I�1�������������H#K��_� ��u���Ay� �K�w��
'�r�l�W�o�R�F{Q��^�)�nl��ڭ�7�n|��v�ȳ���#����e�%g�3E|K�]�חL�������;�� 2<+�犆�r��
�0�B�C��L�H|�u�M��Z��O��gt(�.���ݠ��V�j�N�����b��}��Z�f��B���8�	,������^]�xYY�4�"I#1�(�Ɏ#<0�௉�B:��<�ji�I�����x߅IAxP�Z%�b�[�x�%��y�l.{+���'Ɣ{Cm����wXz`[�d��o%tHr{��a�hXv*�o��I�'+,��$���nafP	B~�<5Z��Ǟ��6~0���8��:��ScӃMCi:*xK���w�������c���Ͷ+b�Ŕ0�Pp-��>AKT���y ��v�o͕8�V���;�BAn���IF���H7
^0��T����H���zJ˘.���|���̑_�W��h�"��b�m��5���KJ���C�f_�6����a'�݅�W��h|!�s��8�,��~���n�ߺ�D׽�!W�Vb���5��]���w��:y��c3.Ku!G���ɂ�\��&?��k�Ӥ�3.��{�r��(�* �7E�UH�UJ<�K`s�sB����:?`�X2A��������k�@r4С�XP�}\�d�*�f /��.�ɠ�j�bsG���>&3�Bf���(�~~����O�E@'Wa/ʸ>�v�Z	�� !f���͋��'���5Nҽ�/�5,��ʄ�rz��]��`����%�b8p�;��[�V���BcbCOܬi�Ps��qs�/rja[qv�	ʊ]����Mg/��iuR`%Z;,��� �f`PΏ{���=�Y1o�b�PXe''�lE���"� ��lX�<8��r��`$���B��C�C|�0ѡ� ���w�`�i�K�B]oeo�.c�䒬n��DU�2A�%��>Jp��F�4�C�eT���+297p;��1 ��}Cb�s}ӁW"x����9kA?X���f�i_:g������
0~#��2px/�鎿sym�fxf7a�8�Ă��7��&敯�#�X^y&�TG��S*wj��dㅞ�i�D�y��u@9!���N�wnZ��Ԏq�W�2	�l�3{��w*/���?�0���� ��	M'��E���8����5+D���R]���=�'��v��G�eFY�NFC�B�(N��t���(_�"��r�>N��֙sB @�4w�X�41���i�����9��H���u������t��&G��Q��rA���[��+����_�=g�<W.s��f:�[s����Fq��M�|D"�D�~�*��"��ot�@�i����fn��o����-I�"�N���)o��X��d�.����͊β*��2Ӏhl)�9#���כ;���'���,)�N2�Hi�Y�R ���ecv�@;�e��\��ߡm��B�"�]����𲙝��Q���̖��u�$���h���Pm���*���>�]<�/��W��S��6`>t�i�F�I�M ���O����ᒢ����H[�ҟ �6�3������#�n��7�"e �2ɕ���3�)��S�Ɵg��+w;�E���T5~rg	~%�8�19�fq�f�M�@�	`6H���G(.�~�x���s�
;��T�5���(9�د�ok?�l�ڹ��2��	ǣdxi,1�'U~��u��mJ��� �	���@�PP`�{�3B%����� ��##�B����]�l��'=�+.S�~wN�0|}�Jt�<u_l)8E&��8x�>�����dX=��6�CpU�сL�u��b�x�\K��*!���D��R��$l]
��@�E�u�L�SD��K��}~��W�,9]n��QX����R�kER�3�4b�d�1{$�Θ�O{9��3)k�c�Ƴ�	g.�b��4��sW-�M�q��f꓄9��N��
h�R��ʁ�hb��,��,E��ۇ��e��Ӎt�ܛ:�jc�I�ž	x�'y�B����$�qd٪���y[��:R'i�(}X��b$���s4�Z�f��tCpZ�a6ɻD���I%��;C��h�������+��`�`�/(!A��#D)��M�tϫ
�PԚ�Ƽ���yp3��P_t��_>3{��s���ǈ�Sv$���\u�J�����g�UE3�$�KQl슦'sж��C]�L� �&���~l�7:4H΂�%�S}j�c�fUP++}8:c��}n@�#��6��v�?zoϏq�l>�����Z湸d�Y^��NNG�oV����2�yL~SL�{uKAL�pe�*�>hl�=�|�p�8
+?�_�4h���y+W�2ݺY���2H�ќ��G{�/9j�XH&�1'���!{ SG5��"�	�Ҁ��d�I8VH�*�������K<�?��cy����0����5����VCG�C<��$V����+�%&�02��E5w&BmWl�u����tmr���3����M�I��b>�s��B�l�3(��|l�:Zᾍ2�T]���
ij��R2�|��x@0���b�\N���+I!��:.>Ԕ�¨7e#tTޓ�WѨ�N��+���0ɤ/�j�۰�(:�FW��m�����s���䃗@ϰ�;co��d$�1�!�p�}�Ct<�P1�2�R��NN乬~!���#l!�(<�^+�$.mC�x"�!�Җ��C�ur��X�yj�!�l�[+��IS�����d���{��M�U���]Ǌ�U���E���چt�Kr�"�f�z�^���¦��r%p�,@���Qb�f�Yպ��0"�<�1La�Fk,����4?�����P�L�7���s$Esg���$��^9�g
V�\��M;r�]9����s����S�:M���e}�ک�IQ̝�p;C
9_Y�-��8����eٿ�V4?PVu��0�a7�$N�k��t�X�"��kki+EhK&��H�-��m+�����6	�S>�(���,�,�S���^��zn��Y`(������;�E7c���|3�lĊK7Ι\|�w�Y�Ċ5S��Q���k�Z��ڲF���{�}�Ȭ[.j��-X��v�55���0�'��xb��~Xm�VD��vFF���mO���]�V�9)�/�PK�5)��|����ZJҴ���V��4�L�F��$�S�Q�
m $:͝.��B��af�yy�9!���v��cG�!naa�Oؤ�H�8�q�
ͯ�*m�+(�$��N'xt�@S߫�5�re?w��DCE�}�D��L��dn�հ�x��S0f�=��?�8����0�����;ߛ�) |�ʟF��*�G�=���
�N'A����g�^R5� ��*Y��z8v"`+������D���f�8�]؅��0NG���ލ͜��}�P��3}�i���a�F&���1�
�f o�m�5�Q�M�^��c<�+�KY�[�ZMfB��J�.��ˎ�F��'��э R;7����,0w�� ��O��ߟ!Ji찏�v�h��k�eJ��g3OwەP��ޚ*�ʧ��p�Nq#<�+���x�,��q{=�]�Y��GS�
��k��v�X�tms�l��C��	D�je�(�}��K�L�K�����
 ��
o<��z��NGie���i�[��q�@���s11J�T��M��#��q�y¶IH�WO���{��qF��6�x�P���K6
��ΗM�[Gűc%W�t��7���!�K(����TD@���#�4:�?미2�= !��=��D�L�����C���@A��U�^F(����|��ڱ'/nFw`�ɬ�
�Bŕ��>�g�~�y�,Zڽ�!�	��1�x�j��/q��7Ë�$L.N	ҧR޼�*�}v��|�ە��N0�n���A%�|ƭ�KI��QI�Ǟ�C���Ұ3�O��#�(�vj�1Z��!2v�s^��/��|�jh�mE��A���scM��%=j�'�+�@ɪ��"����7����U)�D^��?e�+���s}��/Z�q!�����:�<h��v�L^ ̎!�� ��D�rtl��vg��zg�J1$��(��:�p��Ú��5�����n6�F'(U�A]�&8 ӽ�CJ"��;L�m��!�l���J�uI͋��"����kKSq;3]��X"����V$�1����t[��oR
f����[��K��/�}��3����z;��� ^tr�y�,�B9�p_���m�� ww��z��>qY�t���#"^�K���VQ�N���Ԣz���s��\n1����^лt"����R6�NZ���#J ��̹�pZ4�O��� �7�T��}zn����W��ğ�D� �	���{���^'���nۘZ�E`�ڴ1���w�U�7��A5�1X���S�9%��@�'bPp�c�s�+�I��z
����aν
**����2�e"�d�q�s��}W�Y�ӑA��KI,,�H�(���HCP�&��}���r������~��wC�:j8Z�t<$ai?�{�	�eє��V���(��.L�A�I��0���-���"�n��Հ%�x�o�p��Xp��yh\R�o���|��)	�*g+�����ͬ� H�Y��'X��20�yg�i��{�7��g��dj���-�cl��#�D�q�JxA��L8�fT��8ރvw/��׶��E�va�{�9"�֯��� \_��Z��=�`:�V��s�=%'5iJ4O9��w+����yZ0g�.�e�d\R��+�ew��TqK6l��d:P�r��*�w����X^���E@\s�O^p���;�W l�1ِ�b�C��� �2�*}����|��
x4/W�Z`�`�"��+UY�>Ǹhqk�y�S���5SV5��釥qBK��E�i��۫_��F�?�dr���)�M�D���Nñx�l)4�,G�7�n	�(Z�4��z-!'k7V������^|E0ٞ>G$y<C�яe�GY��d֒��L�ʯ�п�Њ0��}q2��ӹ��[{��G��ܜ�����$��F���u�ڊ1��*�`���꒘ �8q��+o�ڔ�_��z<�3z6H�	� ���~.j���W�LZ	�^����,�������<Z櫁^�OZ�� ���zi�I����ݜ��:�r�Z�����##�Ad�˘�>�p��䐌�+0�e�Gh"�N"�+�(��1Vٜgm�}�@"�V�Z�|�=L���'��	�Is�Bo˪;Q�����W��z��L�qe�����+n�UrJC(%�o쨃��5�ݥ�#_��U0f��{��H�~��>�`�(dޅ�0�9�� �_Y4SuoI�Nb�8�!�k<���Pi.�q.Q�Xw$���\�r���u.�Y����0l�`?�d�[���% ���{wz�ݘln�b�ƆƨWx�|��5���3�#DL`�(pE�B<��Y�-��n2������4M�nn���DmbAؙ�Q[y-?�����O��r��B����4�|�hi���q��������S�$i8��f%n\=����L��U�u �n2ЗE��R������P&��,�`{b8X*����e�=,95ɬP�Հ�-H=-�Pd룐�ѫ�~� /K��V���6��|M�$r��xz��}�d�H��p|��|,7��gt��&�R�,S)$t	�Pnp�Y���%S�hG!W�@6%�^q�o�AB�I��dJմ�z��\�qҶ ����T����ˠ�D�G�uC��AI��5�R,۝�m���x�lTV��|��;,U;/E,s�3@�u/;J0�40���LLY0U�	�Ԋ+�r�O�z(<������a�̹�qrD�l�%�`�|�i|��\������s�-�m��+�lS�R~DH(��G ���Z�_�* a��z_FN��>�.�CS���F�z�-�5�Qm�ꓹ	��I�Fp���X2�@�,5'4�G[y'	]"m����g�Y6r� �����=Q�|�~1�1����̟r|��o��0�x�vN����Z0��\8`VË)	�+���A��b�t���w�H�sP�}��W�m؝�;  C���>Z�f�ӧ.Ϡ�P���-/1�&ҵZ\.�Z� p"�������L4�Z���z�8x�-vw�e#�>/�n�xڿ�毦��p��