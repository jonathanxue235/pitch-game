��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C������V����hN=��a���)�硹<H��׮��`̼��D�g�;�mR�#rj��S��k@'�q�/�ha��pc�R�(��g�F�ו�����`d%D��G�qK�DW�+X���iv�O�O����9�t�0���`�<�F�2MGJ�g_Ю3����Na/��4-^}��ru1������>�9�Z��_1��uC�wx�cn�͔�*�������P�v�,\���)෾�3�n~�2��(��ȱł�7���!٭�4�3	[	:Q�ݡ*���y):�:~Hm���]�:.��/��@��(��<{��ֵG
�k�_�.�װB�'C��B�bf�i�ޅo*(��k8O��z�1��5B.�B�b�W����9��N�����z�rvc�pr����۬9�"źN�pȇ��K_�
�G�m`�ϼ?`�$^�61R�D���+��0�.g�O�c�~J����r���D4z<�y�'�
׆���`�vk��fv�H�p�������\L��S�%��7�����gʂ;��H^��o{tТ��{5�P�o/��P*<f��̧�ъ/��N�rI�)���|���U'L�Ԑ�X����k��rt7�z@E�0����*-��Ѱo�f�Z�To��l���,�	���b>P�&�����>�5g�#��ܜ@L�����eN�J����k���f�e���F��-2��_�%�[�h��O�_Tt]�6j���Z�����UT_��D�<^0��S���AG����f�Y沩�8�8Jp�활I����J�4�I�1���1(L1r�{��O�����$z?W��ܘ6�O�m�V��"�n9���43�<������c5��g0�>z���н�uq���0P��Ag��V��a�m�=o�*HN���!��)����珱-�tS2��B<b��40��
K�U�ر�Cr����l��c��9���p� �����զ�FnƗRl7�Hdh<T�;`C5	͎�z�oC����3-d�Q��L,J�	�+��8>�����=� ���!��b� o�\�_�DZ*�T¶e^�Kh6But���t���L��}M������v<;(���
?D���1̸�෺0(�Vfq��O)F����k2y{`�1�E���t���M.>j�jx�J�@[a��tI� :+�N���=���Ě�<��?'܄Y����0H��ώs+<��M�p�Ku�v�o��
3Wa,/7q(��#2r�U`rq>�m�j�������w�m�Klƫ���.U�}�1�}��(��1q��%JIW��)��m�m�8�64Pm�=LbM��_oHI�������	d�O�ѷ���m�����IqRO�����P.�{�X����!��R[2�9���)ё�I\��Y�����Ԅ���<�gM	S�(]�#�@L��!3�JW���9��[�i��n�ZmY�Ń)���tZ��i�o�uث�}�������B��֩"D�[/?b�4�_TV�´a�P�OIF p���׽�J� xH0�w��@��-#|Q���Wf~�-�H��k�@��[����x7� s�v�;���lۖns_�k�j#�{���" ��mc��Ԥ�-��S�3Q[��ĉ,�� E�,��TN�C�Nn��9��p�j�k�w~B��ыI*^�D%#����4}�M%�UT5���5�DB�Êȷ�;��]͹���d(���d���(<��������0\��e~]���skxv_��]h���
HGk�'��-I�Ue�\ėuiNBp�9$�ȇp�dd�ۥ�4���N��7������f��)�m�(^+;B��yI>��T|Y{_xwm����f�
v�G���D���R2pY�I���<P��86�i�]��L��:���+X9���3�E��Q�'{����*�(�H��7��!d��N�}��U#0�MI�(�,D|��ρ�A!o�F��O���1w��|�"v_GK�6<X���d�Ɏ�F��G]*ȶ���&��D��v
F���_rtnӇ��K�8Q����l�@�J�<q2�eV9xy��Vȍ���=:Z��[2]K�����G<y�K�zHRuW�u�Q�痤��Jw���:)%66!+����B\�wi^��T�Oi���I�cK�R�� W�I#��Mj �ty�\,���M�I�#�o�.΄���j�3h��f*��b��u���J�(T��� �ڹ!�f��X�	nU����Rg]'1�a�Z���v�eKx���v�%s=��^�����ͨF�o��i(}#|(%�P�,�5g7=���wy.�uOSC9f��0��1v_.��sZ��ȁ¶Xf!�5�N��y���������ґQ�� �nW��yE����y���%�.jѸPx}*Lw`5