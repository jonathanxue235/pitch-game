��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� ϲ���4cg�b8r?��F���J�f����@-�$�;�R���\zaQ�8u�%�l��e�1���W���4(�Im�;-WA9_L��g�t]��c#]ژ1[[�:��`(��<��G����0z�a�I��B/�5xb�/{��#7����d�>!
Q�bc�ӊi���0�sF���hwNK��+^���"SO�^��Xu�wxKHI>e���:�8���J4��=@��eR(�6��_gx��c-��ͷ��9([.���}/Dg��8�7��S`؝F:(�.��Ϡ�6$~r�Zw��}�١�J辰u�
��9<AH�{T��v �j֋4��
6e�s�g��`��������Q�yX�y�'����F˒� �kGx�r���'T�u4�6|]g�I�����=w�~83+�#+��`�ͭ�Aʣ`�ږ��zt�zfiy��?-n�:S3.�^[}}�o#�D��s��⢜�z"2i��ܗ�W�?������C�j�	X���%�	w�;��G�.�b�]�>eb�e�|#>�9F�K�{�V�2��h��!go[ׇflX�X�ş��3�c�=��	��O`G�HWW�%�1�ݰ�p����6cY�¦���2>�)�-�4��:[�#���iKfVm6_���C3H,��pz��O��#;|ls�aۀC��W�%���q���o�?�#֟��*!�~Mds7�g��N�±�Xg~G��d�F�hx�C��ä��p-�S2}C���7j���Eb�Q��gQ� Q ��������˻X�"��ű��\t���@���痄[w�l��>�\�_�w�W����K,��r;���Q<#([ۂqRs�_��7+��b%�(D�PUL�++�(��Ow�Ö"��A��!��]��\�q�t���y��]�ȾuT����)�;��g�*�`@K5��瀲�io�@$��d�m��q�-G���Su׬.�,�	!v��xeB�ʽ�XO�ׅ!!y�7�Z̘�A'���%X� /�)��)0��"��+?�*����!3�! �"�����a�'�����|"z��'v����욤�:�e��8�&��s��書9�8��b9ƽ������W�k�m�}����	e�����!��W��O����h/��y}�'&&��r�FAh�2�{\����%$��Z�r@1(7�x���K������{�E�j�l+r���;���8p�E��O>/�=$������˞Ż�A��>؈�8�U(1�of��2@�x'Q��G$�i=�v�Uƀ�1���L[�"9J��yyz�HιM9n�/;�o=�ߚF@Xa9CᾝM3���=���LuS�zd�YUԉ� ���:�08G���nH,:��U纜v���Vȶ�1�n��A;`'6̛'�ʓkDNn��������F�7�*:!����(�~(�ZP�"���;R�QU'=��D��b�N1���J���ڶ�5�v���b��:�_;mpa50�t�X�A?<Ro0_E�SD�{@�Ǳ�e���t%T_�5��0������!s�d&�04y�H�/�m�Hz�&(�]c7ʪ4�=��m%�?q:�E`ֱ�¼!�&Ja�=��;ɄUn�k�b�p1� ��?�}�\Z�V+��ɺF�tQIW�TP�3��W����#7��RJE����x�,-���V�����3Ca
��R̦�P�����J ��s����',�i����1�r����F�ȰZs�.����ux������jc���i.�QQ�#
�n"n�t�/9-M��<��g�&b:�o7�s����lJ�oR`����l�1y��b��١Y�L��������P��������_�ZUv�C%�Z��MDG����N�=(���И ���oOf�@p`6�IRYǚ	�40��o���ش��dO�ꞛ�2ꧦ&m:�{��1	e ��iF�A��@����=s�Tm�k�mU���R�4�V]2�v����B�_٥=�#'�����ik��h%=�����1�����o�2���jt�S�/����_������pҰ��������?�$�����жh>�̂����3�↥cjC��4��N�K+�b@�s3�]-ȣ�����+p��?��ͽR?��u�v}�#	��01G�41\F( aa���w-C�п{��"p^"��P��!мZ|R�$�$�[�r3Y�o���{��ǾS���^�t�i��R������W���TqlV�?�1k�ZnOs<�kIu�PJ��O����p�:����Bbpq�WYdh;�*f3=�S�0rP�I�=tp��-��¢wn��p��O���#�t�[u�H�o�ڬ��+��2I5�������nط����L��)h�.���i�<���D ��1��Sqb���n��$'����r)�
z�l5k d�db��~�&d˼�g~Z�Gd�U#S׃��%��{�p{O����z<�c�0�%�E(���\Wx�a�|�'a��[�
�:u ԉ	��..�Y�E�g��J2ܮ��C|E��x�dw��:�1����RE��.9l{�ނΨ���q"O��q�B��$��X��;/V"H���C�j��P�#pu��
�ŤE��*o?��ԕ\�:�C�l�
�R�Z�/u��f��M�H-jZM����-����,b.'�0�N]�s�;ƿ����U��*T}�r�I�UBp9�F�;! K�SF�,�5�!���
�S�bۃ:�n%�h}9�#�^1�Ј��2�"��m�Z���~���P�.NvFv���l`�Sq{r����&��4D�lL���9I��]�L��^\H��M!��I����%AuD���H����
+j׽���Xמ�(���j�bQX��I�`v&�~,G^άkJZ�~�j�9�  Z�f���˝S>�����/�K0�ۯ��z�^�{��Z���"ʡ$�;�����Ni� ^�3�8X�Z��^�le���::��)炬R���{kktCu,�.����g�f�C��m,�LAK;�L���B[��T��{~qrb<R�p��l��"���N117t��]:f6+�*%��jג$���|�5��'��(��&-��	p�㺥kr�r~>�#Cb�-�~z�lFe0s%Rqà���1��%���!�Ez f�N1�y�|p`z�0�d�a	D=�D&�A!Y���Qj�Zj�E����(n��4��]@�G�����a(�L���6Ӗ~9�U�_g@cRQhZ�7�}�a7�ް�Խ�����@�o`y��C�y����*����A<o�F��F���c�U�9�P������ߤ^1�b.��[C�TMٞ�K�[��՘��w;D���-z�>��ʃTj���Kg
���wE鿅"d �w�c�WnS��}������F薹���?�Ia�G��
`��l��c[T�q���gO� ʻk��[�vcj8'�^�n���#�>�wj^Kʣ߀�+o�^ 0��o"��������(�~�����G!�T��O�R��#��k=`������5��D�S>�x3�f��� �,�f�`0��/���L���Z���HHن�#�YE�\�=G��ct�D��(��{�nΟ�?�}�3-��w&+9���r���z(���=_0��F� Y�Y�[`@�eMY���Gw�W0�ߟAK�Y�c�����ؾ����Ef�۱�� ё��ˮq�c�>V�X�;�yp9F0W�uU��B��ʶ��!�8gC;��uc��<(��n�r,Q��n�
���&����Փ[j!O������6�}���X>����@�$K4����� ֳ}XR��)��G(��=ꞣ������Q՚y\1�C�U�XK���>ѱ���I�]��Š���$|�L�J��Ϋ�씄"�S���@�	�x���޲�}r�G��[�f�=d��3����y#Z�'/��9�2�FJ-	��H��\�zŴ�^<�_��5XU,�$������ ��e���#����l�2��`r�3B�cz%>8�梫&��n���]�6Ɗ���t�%�����֙�����`��V��!ʉ�$9ma�����8��� J�4�7��b,�T�j�v<�.���=£1ߜ�#�am�0��MћM��
ٙT��u�ƘkW����H1��@i���Xz3�iL #� ��hЀ�Y�� �Y��x%&A���ٖ~f6񣝓,!���j���t�7����.ǥ��o�{v��Z��~��ß���&��]?�:�f�ɡF���pv��ۨCm�p����K4��6m/7�<�w�򨣦�E�^��yR���іs�@KP\W�_c�M}�ѽ ����ܱ���0R:���RN�6\Q��c�^�Θw]Ȅu�R��o8�!:�� 6;O��h����>a$CoM��0�w�ZH�����n��!Pd�1��#N���}��K, x`<�>tk5z�Ψ�Z����EJ�8����'�N4��'�8��֠jQO.r+��M6m�2�LC�� �;�p>"�g�hI�7T�95�;O�u��O�Q����B%F���`��m$ޠ��l\�%���Q�KEֳ�W�o���ATd`��2��ƈ�E�ڍ �hL	x�ơ(��9���h{8���2���'��ԝ{�~�HZs�@�T�`�x��вT{Zs\�1��r_���O={n3��J[翁u��e�q̉li���4��f��YېB�|O[ԭQz�t:轏�ʰ��Љ�����+��3��)���.��A��4�%B��'��ݚ���yS{��@��|	�@q|�d���q�W=`�˒�]���@�X�s����By���Zj���^�dO��tl���(�"��QɿЖ0E�>r���+x�s,�Y��2�0dZ;����Y�G�@�[�o!��rEK~�O�ߴ��	l7w_#RU��A��bJQs���[�����e9վ3�q>��v�� �17�:<�8K�mĔ�~��_:Q	�Q�	3[l�!�M[�Nӆ���KT�3&�JbH����;A�=5��J?����C����C�!�w�rE��Lp蠸.��{�?�P��j w,�V)1��M��Mcm-��O�{��׬,!�~�e̓����ˀ\��L}����ZQ��#?���D��X0��������V���㾻�dQ oc3�=�zxs��Fz�������-8��<,w�G�]�H���{�������e�ы�})� "WI\>#�;R�|�bx��-WS��iP*X��_�i��?Q&��@F�B74(�X��̭��Y ������fZ��g,���R-HO�<��G�X����Cw��bt��7���2�jϛ[web�sƼ�oB3@��a���P��ʹ0Hظ�ظNn0	��]�}�Y���r�w��R Sr�����Rn��]s�/�i�=�:�,%LݷQ�X�FP��o�l$9�M�3޶���tjTZI'&H��_9{���f���l�C��%�
���J�+A�R	o�Vw}�3������=a�g1��-���b�h���aM��_��:To4V>�?����/T����d���ë�]��+-���&֬�G�k������ۖ��O:�E��(>�k�1��&=���}��s���#��tr�B\���l���Z�����B	bY�9�.�t��XX��
�����$��T�_+�]"a�K<Ԡc� <P]S^��\���E{��*�����~Fq`��2{��W����7�C{�y�W���I��b`�k����/"�X���s�Ul�����E��Z�U�9�Ծ�������/o9c�!���S����B����@��Dg�m-3�گf��R/�x0:9�2u��*�H�&�y"����BEvPc�="a���K����(nKXe�� ��f_zv���[